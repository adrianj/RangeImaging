��/  �Xt�`$�����My<~}�A��5@%z7�FH\�0��-�9EMx*1�s���v�G���n�2uO#)�Y>�P[!W�n)6����o�hY[�ܾʰ��)�q�3����ϺeK�^)p��Hz�{%,rU���_��^�^ۜ���l��1An"3�"�����o��LV�laD=tp8FΡ��'�N$4b<9^���_.x.�S�}��_�wd�rV9Mz	kb�X]!��:J�#�7�{r��x���:ό���Ȱ�2y/r��m�\�R$�<�V�1Y ��\?;W^|�bAj������h�W<j4�U�e�c�ދ�c�k�1�xix�`J�_f�2�	�ӊ�Y�������-�#����R�9]#�G�QӠ��
�N�< ��/F�+*��?<��i�/����b���X*�ꂖ���c �c����Ҭ�rsoEAC�XZ�M[��������}21�N/'S�2��b� eM�x��44�hVk�
����*6	���ҡ���㛜�
��>�VCޗ��9@�ܴM~�����~���:�[>�!����W	)T�F³�.�sA�Z��R�a����F��S:YB0:�;��Ť��27Xaϙ*);���%r�(!d5cbj�!/Tל'�N�!�w5��f�_ࢇHڊ�U���W�q��)����b"���bM��T��m����7~�.�<!�o�0��`�ˎT�˼�c���&��;��Ў��<���ƞ��s��X�r�Y�����/a>��_�w����9i�#\����h�c0�b�\]Θ�%`�@] �:s���m�d��Z�s����F�f͜��p&GqC����ι�L|�P^L�&!Aw��x�9U\�+�f;�jI�(��� 4W9Lru?�F��'a������N~���B@M��bf�9I"ei�j�ySe��r�o��g��qP��&p��M�����(qK����4;B�y�>׮��f}T�"�|��f�
G��՗$��`p��Z.��T�F\4��hD���x��O������ū��D�'�N(cQR@M����饷���a&��3����~�~V]�"N����{O.���ת<}�pgU��Y[bЍϠ�g�_�̿��&�WA��܄�Rv���c� ���0t֛ӄ@��2ʅ1�AR�t�@�g�,dP�w-�"����5� ŷ�u ��ш�AF�|�:(�T�{�P/	��a����VJ몢n❬�_d�3� F��x��0�b3� r�q�]"lΰ�����'�����1��������Q��X�BY}�+�����n��1�z��aR��C3�o�l��(~�ߙy�9^H��Hĭ�[��m}옳�+=J���J�U|7�š$��.Ԛ0���ɜj@C��T�l�NQvRo�v��]/?��\��r�`�:N�$���A*͏pa�k�����W������9ӜR,����[�7���A�l�����E��Gu�Ihy����fuͩL|���B<G�����7��Vw?i��n ��L/�Ho5#�SgRo�
`R�2�,4���JT��|:F��d���F��y�^�N|�y�3Y2�,���	��M�W*4�޹o����;���A�$9c7�B�'!�ךּ�h���!����F�T������]��N��h�n�� �i��J ��Eu�f�o�h	<����K�q�hp��K�:����A9M�t[�����bO6ܾ�
r���#�+�s��S�L�H�σ�����>���m�rv%�בo��9@<����MZ�U�V�o)�&hh�n��3:Z�БsKC�q� 8o�~�$�2��#skE4��*�9��dךgH����m��n��gZ��)��L��WMy�4�+���CI�����W�$<�4f{���$-��z~#)ٰ��r�ɒ��z>C����'��4=�)�J��Ȩ��IY�̯�
��~�)Y#��`�I`��A<�ii�r/�p"7B��3s������*�h?�B+��?�d$Ƕ�(E�N<� �]��x|� �Wg�y��9zM~��#�W9q�?o��	[�i��_?|G�>x��ۚ 7�z2��sô��^\�{�A�ˢCB�������@�b�g�q�6����ٔA� �1��"O�y�V���L*�H�C��	��Mx{�5yc��;��<;���� �F;�]��n�H��WvR��VFgn��f|��_<޺`G�i��x�@�ou��/��F���N�%1��J�È�@SN���sp�$���Fk����I�ǃHF3	��A�W1�b���)��v�[RHo�[���g���~f56�k-Va��VH��^7�+���aIW�~���k��JԀ+�<�`��B^\7�q��R���R��EA�ǈ����s�q �9��E�[BN2��LdR'�fa�)~fB�7919�e���{O4��Ӧ����*<0l�sߡ�k)��g�ڼ�a>v���	��3�$��\��i�����N���v=����g�?3�E�ې�C�����2%�y���P�� �g��pq �pw��F$T���RμY����9�$�V���7�+}*��sa��F���O4�Aτ�Bjؼ<�g_)��_S��
�b:�l��u�~�y�/F��B�.$�t��紙P�~ I�IWm7�m�6�Zmve��B�[i�.���!��	�ɦ�?�I�$1����N�R���l�͇j��P�  l��+6���8E)��"F.6�Ҳ?�d:Wt�&
�C�#ف�}�i&�i��Y-@��#O�`��f䟣ʾ��wN�>��CN�Q+�oة2���ܴ��&�� K�og�!~FaX�撃wx����.eJ3����:�q�xL,KG��/�:�ũ�r�`<`s� ���mADvh �v���^������O3��������i�j��\��k��oɓ�|�'P/�W7���J�%�;�vD)Q�[��u�F�seb�-S�&���H���j�n	���ˤ��<nZt�Z����~�(?�m���{� 
3�U��"o�<[��y��~��k�4�B���� չ�LsDs�z��Ӎj�گ��Ў��&��n�v�г�lk���%H����D���O3�2l8�y�wQ��7s���X*&�f-Dn�&Z j�/� h�z�?��-4�K�<�8��I ��s����3���d�qu��p�C/���N�����S��݀YZ�`���D����V���{�u���A�̱q|�j�'H3jwȏ�Z��1��h�O|�w,b�P\
��!���6��-t�L��X~3��0�G8�����n��N�xEq�eNհ����h�!��a�ܕ�9����x�6�-"~���3-J�2p��T��O��Q)鮴i�	�+�NK��|���
Y& �d�R9�+ٮ��=ޏ�G6T�5��=�Yڻ��0�m(�H/�����@��8�q_7-�(��H���w����(?���R��#	M�K��%�U�p3�ˤ��b񇐆}��������TQPQ��L��nl]H-�0�_o\?8s���Z%�����a��2.]H�r���6��t_
������ɡ5�,��&[d$��wO������r2s�.��P�"�!���J� [8E��s��8Bj�sZ�K~,W��!����HׯY��G���iK����oA�#�)Y���C�L�j3��^"���b�`��s�<]w�JH/�4��s�^g �G��{4|;��BVb����ld��D%h��~Y��罢�����S�I4��B�����\�*����+6,x�=,	�����!L�qrxJCr ��g�s�"���H����-i9�~�@-�t��<�L�G߃��������\?Ƀ�p��.[��O	����Q�V�ƒ�h[ː�����D��2Y͈�� ��z��0��[�d5�R*1H�Ŷ#&�����6�P/~@/H'��^E��4�FF0V��T2��P�$>�y��4�l����o{X��E�����AƆ��J<Jx��<Đ���2�w��D��6��)�d.X.�'��k9���n�8�e^$��H7�w��~�&��]���4�_�CG�a��zpԈ�#Ew�F�浪唷b��o���5��|з2�Uԅ�%�T:ՙ�z0G��}e����O�;�IC�����F� 6{�xB�6��gf$�W�ڗ ���U�U��"!�Ous�\�Ik
����S�:�󍘃_o����rG@���tP��-���Ibo<���m��.(���%ӗ������=��'p0*�����sœZ� {
���w�g��,�,��y<�Q��W��w�.��U�V*�A@�!�ǋQ"u6d�dG0U�޾O��S����S|:l}��R'��
���r��6��î��b�3���Qj��ݖ)� )Ӆ��,3��\�[96$/�J�]���Y�Ș���f��+�p�N�n�+ŉޡ]W��ԛgR3���[�3sd����9붙��"��m�7r���f�ɧ�:�`�ZB+l�5=�ѧ�@�U�VZ�j�v�d�_Y��2B�ÐI��`������F����#Oq+�5���,ףb����(�լ/����ѥ���Ҫ�����)?����wVj˒3+~�����V�3_�ӓ�ü�Z5�ƺ������%c%,�E��C�z-���>_�'m%���owu�����|I������~H�(zQ�d�Z�>�`	��j{ҡP8-UP4���z���s^�}%�l����$b�������!m��#Ti�v�}e�ҐQ�م��%�0�|	)�&��(��F~�5�w:�N&��d�OJAi-Wwk��LC*�QW[t���KR�*4��ȓF���F�,I��+�
��5O�_u�CSZ͆,�+׸����$-�QLF6&hS�ׁ����&>l�]�J|.�,�P���ˏ�T��vP]��Ƨ�%������GQ!5�U� a�7rQUM`oc���
0����^Z��P,sAu_�E��7��0�	��٠}�w�7��~UL��f�R������"�Նx0�XN�nfr()�<���Y�1 ��YI�O��d?�ٶ���-.�[�9Sr�^l�y�F��.�O#64�қ�0�)�dIYv@�oiE��Dy���zWq�y���w��B'>tR�� V�G)m��M�E��UB�t0��D��]q�zCA6u�-�0����~���XB� ''���K	&C�?�׏1X!� |{-�Ú�ك��8��;0=I�Y�~cw z]�oZe����S>L+a�<�	%]N,h�Cc|�P���z�V�3�K���j�<]Z��L�lBB_5�cՈҮ�Q7D>�RLN}<\�,�]�X���խf�s�����1L��G���A�v0����o̙����d��� Go%�3���V�҂;��rN�l!J�#bia��ØO1r���.�[��_Xc�Iqh��U�۳��_tnY�Y�GCq�<�l��5�'�js:��٧"΂;���<��mni#h2�����E�v�T�D�$!�'*��p���p �(N,�:9�A�4P�g��B��Sβ�*������۩�� Ȍ�\�u*Nb5���a��&Ʉ�<�����3-td j
��_����<;Ђ u��n�G��w�\�FR ��������������n.Ca��<�>w:A8h2�Yi��޾º[h���z��h ��&w��lb\l�"�a^tD��(��O@D�=棘�E"K��,�����D��w˻J��V�yTS��f���`d�/��H��=�`�����s\���?���+��>aB	�'e��ց����̫;�_9�| ��`���Q�NWt����/�q��z���]��`_�qA��4ƥ6�g����SXA[�ww-3(.�Q;q)�����M<4����Z�>����Ұ-,QK�1�l���$���v�%�̜ͥ�%�K�t�;Pꎆ��|T��� ��0Wj�Ib�������_��V�U����g-��th6a���+H#����<�ihz�� ��5��D&���� �����ћ\�0���{=��bH`�����̡1�5T����{���o� �������d���1� V��b���\� #Ɩ�-ܗE��x���\��1��si�\m�ٖ��T����O���A�Z$j-.�p�	��g�®�>�V*�[��<-z�(��ü]���OX�d�i���?�rp������4c�f��硳�Ǚ}��^L�_,�]u��w�6hF[ץ��*V��y�
�����:lѲ�<0q�Z]�'8����n<�-�ϐ0��ƠV��T���QD���M o��b�\4���RK�94���]����d���euA��|�Chv�+�P�:C�_U�gkb����6> 5T�y4�����T/�̝�;V�X�Us�p�7��I���24I!P����;�r���ŝl��j�m�p$o�[5�95�3�F�|�qu�v�x��Vn�V�|S2�V\Fif���?a�T�k���帐n8פ�h��&�JisO ������6n@<�����-b^x�(�	3~r�(��u���l���"�߯�KY�t����(���A�n-{x-`���p�_d���j
���z<�y˟��tP��]h%����=o_� <N��/�R��GZ��}�0��[�\��ҁ1`5])N>��8��j�`ɁS�aR�rlL1]������;Q�P�L��E�m0'
Ԍ8�	��q�š��4|����b���e�&Rv��X�n��k���zO7��@�.Dr�(��Hyy=يEk�����+`F���Q���&>��UJ���QYcP�2������AJ�E`�d^g<>�w̼ugƢٜ����tpXhW��Q�Ֆ�l~�@�ky���o*��� O���v����F)�p^H��A���z�'��F�n U��|"G�5:������$n���!���@s����C��8X�\ʹ\j_�In��ԃ�kx[B9�D�?+������ï�~��,�k���l��껴8�K,_5�y	����^Bka{ڴo���Y: �ՠ��*�'yb�v���!�g{^~��nk���fO��%��e7x�48ߒ�L�8k�`3�a��H���\z%���mT7T��I�ܟ=3�+��ת2�R-�1�>z�f}�+���v����E�m�ZKjӳ���t.�bm��l�����RI��\d��ģ���>/!#�K��E%������1��]�r8��:�wM�XGT��:̯���p�%K�|�Qr�&*��� U4�"�m�W���������(I�T���H/���-��zҝ1V_���>��u���[GGWK����O� JT[>\�m��씧�4I�:ck�а������?4qzQ�dU��fF6~D��\� =������?>ra,N�o	�姄1a�\:8R(G	�fZ�p�v��)���"M���{JDm�k�rm?M���Y�'E�?�~F�{���2�Ƹ��F�9+��7�]M�/�˓`��lǗ��2�G�l�O�	���<�U��r\T�p�&4[p�O�J����4�h����w�h����"q���H� ?`<�Z�y���ӐA�|��cX�V+kl/����	�R����"7"ς��P�r�=8�\�%�5*?�^��ȕa�0\i����`L���=-	+@ ö�KB���w��/��h)�e<ܡ8pcs�$�Az�vB�� �ݱ%?{ꮃ�M(jI9���*?�L���R�Q!|K��o4?�V��L�AK�fT�*z���F=р�ҹ݉�-d�<;�f�[.x~ߖr��E6�;řt[��Kԃ�Zu�К�nV�J�R��,.����C������8��a{K�?����#,c\2`{xi\̲�n �劚����U~�����qh�ݤ�8�!՜�0�FPė?e���^��E�#������/�l��� t��Q���i�,���F (eD����g���Pk)�\&u��۸"��@�aba��� L�ʥ�ALa	��Ogn��#r�$2c���[�6��@��V���^����m(�T��7�约��~1F��K�
�N��(���j(CJ��b�.�YB��u/��Q�-�%��g<�A��z[Dz[  6* ��E�5��t��ʾ�jX�503րm����k
�����#���H{���n�$�����tQAg�G���}�9�d���a�C�'�Q
&)S�zi.#��#�w`�&2��Oϩ-���hD4�4�f0T�a�J"���jЮF[s2ޅDq)e�-�}e
a�/D0��F<�F��~j�}:�=X��͵�a�U��W�)!
��$��;�c&ñ6���{n��c1;�	ҭHH셰/ـ��Q��o�H �n��]W�JM�h�^�]��l��Ф����b���jx�!��P�����/)�����)֒h*�?
�Z�=�z̛�X��B&��m,��W��O��f�; ��g�~�����?|��8�?�JNj��T�����mVN��E���b�xQ=���]3-�����u�`p�V�.o|���	�̮���.D����Mp��"4�ZA?s�P����{���� +�(����0$�eYz�&�\���kO�#��ϝ�dǀ�}�$�+9i:��;���W�퇋���+��/��Q��Z,D6#�Y_!�tlLGK��\G%��EE�+�[=m��D�����1|�]ӭ�(}OF� gW�B�����6�\�8��zw��{��ʂʹ�^����ַ����9�I6u|o�E�y.��矈��Ink��������<�����-��:��T�56PD֐/z�'OR��V�`�3>��>�e�a���
A/^^���m{ō�`��ι�y�a��h��0j`�1ǈ�����K�y�}����x��m�@0�#���k���j ��;�ׁ�l�)�,�/�y`di���3(�(�����_S�y�v��\W�	"�j�E�o�&������oE� ���b�fѧԳ.��L�������9گ�ˑ�UO�T�^�2��7���8�~�7d���e��5y�� �dΈ����]]D�l 9��	5�ZL���J�x�{�͖�${!� ��(������RnD?�A�D�#M�n�Q���I�qg���B��ؠ�'��G���?��B�A�;k����pbF���py��mT��e��S�9
Ouw��]����ԙ��]�v:r7s	��6��w�V�G�����<	�_�()V	���~��zF5O�U�~�;�رXҮ��`ȏ�;K�D�YHz^�9��ub���bs�ͥ�?��5g��i�`Xa����8��RoFd�4�}�ɀ���@�ϦAd���;�=�.�Ny�n�U���z�խ N������iD�m�"#h��Ctc�t�2o�k��WT��8�G�;�p&5x����yTua@<H}X���a[���Y�2���G̩���1�~��lD�v�#�WĀ���iI������ҩN1���D�R�x�!ջ��sfM?T�7��78\��X���8A/u�0�V�_�Ls�=O�j�⺿���d��:�o�V�f����c����*��)h�5�-]F���@A��b���g�Xj3��r�Y7F6\� �(Cyg����c����[���a�R���yA|�#�`��t$J�KZ���<�-���>��GIL��?ݘH��IQ��\Y��Y�+�wW�W��Y���,z��)W�ăM8E�V�������6�#18��@��*��{�����>賯���Ɯ�d��*�p�!6z|�{X����6a B�n1�5x�p�B=�Bn���/sTPY���`J�S�!⥂|�E]��4}�>���S����K�*E,ΐ�G�e���=3$C��~XkBKe:�z㓳�)�����"�^�}�T��%��&>��P&j㇊Ű�g�.Q��j)�{	���U.��P%���R ��	k�Ҫ¯ |�>o`�������]�)�6��(O�:��9$��Ȓk���Qt�a�G���r|y�n�g�2�(�.C9u�O ��!���zYLק��z���ђ�4c/����j�q:R蓧�d�+��x��2"	Z魴S�[�	�e1�"9<
��ķ0�����3X��5׹T(	2��c��J�&.��­gʠ�٘� w�3f�g���|�1_ s
����T���(ٞ]�#b�?o�މ���[�
�SԆ���@@?��JCR�ߋS��_!�oU���+i�)JK)*�op�0��N$���>o�(C �̂���	�� ���dX�I�,'b�M�]Ţ�Ui_M{]b�� \��FB�rz��3��B�����4н$��!��,�ʜ��8nG�{H�޸�*B�W��5~�`�Z��Ch�_U�����	#��j_g�0y�Wi��cVCy���p�L;�l�x,P�M)6�ܳ)��S��a]�Z�1�Q�r�NS3��Ǻ�+���8���3u^���j���q���7�d%S�3���Q�d�9�T��������8� ��3�4ޡ,s�  6�S���LAݚ�wO��:y�)'#�̆i{ ��p2��xc78�f��)�c�q�3HS+�����Bޢ���	a[�R����(��.ֵ�5�?�'����7���b}��yޛ,��Z��g�|g��\�S�� ��!X�D��p��$^�="]�}��wuP/7\�ښ�$ڰ4'*�@v�/t��  ^+�C6�jHC���/���u����2J�[]���׳�`m��9���8�Y 5'*g<��荞K�XǛ%��y��Đ�� �mۗ�,<��`��):�[�T�Q�^�����vۅ�p�v��7x�^�u�70!~�5�5��D��k��m}�޴��1E�s,��u���]l��M�<hM�|��uF�"�s��
h��;��v<����ed�$�T�r��m�t]|�6L��3�q<����4��*��N�Ŏ�@�X��Ã�/�; �m]�V/�H[����إ&%���U�h)��2б�$�^���"?�C�^�7���`/x��)���t���H���r���O�!|P�Ｔ��g[�ӿ]��9�o<W�k��^naSԍ�ǾܽQk��J.�ڵ�o����չI�E�S�/�&�D���^1�O�Q���H��S�u�H���Y�����l���Z�(i&����M�k	3^�����,�z�7Q�e�&�{'/V��r�,y�����pl��/��EE~���H8�<��[�έd7���K�1��p���	�� �s@ J�/�A�֚��6�pS;µ� `m;�
��p���\0�
qVxS�E�sy��P�o��f|���u.��5�"+�{8hR�����+�h����Ǝ{�5��P��B9�b��s֌���!�	��S�F%��N���ߣ��lu\"�U4�����4xy� ����?;�=����\�"֬�s��ґ{��dFk)N'�ז:��uķ>ɷ|����L��In���~�=>=� g�ޥ��]�y�&9��Me �7�=���~2��#���K�Gj�|�/,�����/~���&�|��g<$��E3R����Տa�V�n<-zE�&L��b�L��/�n(A�4�߸@|��F�����`B�����<�N�[��_q�h��,
�t]��ky�;�/�������ԋ��ê���/	�oMg�����=6����+ۻ' B��Վ�^P�(=s�0������-ǈ��|��*l�*��N���p��5��a�g���lR��8h���M0�$فLt�M�]��F�	��uzu�M��|9b����fkn���?uF��I4?����PٚG��6��>��b�u �^Lgk��d���:2*���.��4�Sf���5�x!Ńe4��aؒl
7��U�}�!4D��r�����=9�u����b+gFhJ�i���(����� � Pm������MŻ�w��D��ϒ�n!^�8^��+���$��΃^���U��Bh4%��~,��{5�����c�����:��N�c#��)Ji6vC�K}?�,�����-'�
�R�:9�*8�E����i��E�w_��#�H����� (\		�����uoKC�^Ae�@��RB����R��=� ���L�P��� ��ܦ'N�U�Ƕ���v.	^߃8�a�G�/��B 9� �EbE+δ��9�pp��{������S2�[J�Mu�����|��6��W��W �u�}��[��qgE�_�KM�k�Z�aG��B]vpm
��n�6XRH�\����i�~7���"3�v�}Ww��3��0NW�0
�ޡ��"�RK��W�ĎkҀ�vO�f������yx���kL���t��v��"hl����8/Tũ�Z{��|�H!�D	���'�e�G�=ˎ�ǆdD{E�}y��4�\��'��v�f����Ōh_��"�� F�;X��g쫪�����g���O�e���m����.�%����������=74pd�Ӓ_Gӓ3p�K���P(���lZ6�2�[t�����8�I8��a,eC�7�����������,��3��=b,C��)�Z4)*mx}0��}'��Ẁ��~@��.���y�������R	{���m�O,�����P�/�ސ<��G77���h���8>���E�W?��sH��Z�H�L�dO����X�o&@��a�YT�J����5T�>q���%�'�ƻ�yT�B[��^���U�����!�*�'<����e��]S[\X�&��єI�RHU��{���Żb)P!���6�ߠB�������*1�֒9A�6��R}X^�5�P]NF�e��Sv�8��ܦ@9���/]KO�����e����nld���E7c�����-��&ܟ�4父�k�~6��Q���O:�ߋIj���{��M�YUb�e	a���3T����	6��`�^`��G�|��RQ�Kɓ�
�y�)
4*�ѝ!"�&�v� �������D>��"P��P~���F֪�Gk�+����S���%�b�T�$]/����1~.�1z1	,����K��\+��ɀE�/���8�G�lCHN9�m`<�s{gM��g��6�n�|/UI��kFg<�o.'�י���rm�/�/?�� fM+^� �|�2c�5�%�f���Xl�q�������k�{$��({�+N��R�����YHe �:�d�x��vh5J2�-��f(gB	�ِF�>���������0:���]�|ld9����l�8�Q�=��G{#X)�/��TJ�M���}��{�Qf�CCX3���S�VI�� ����Ey����A�N����=�4k�@�ʛ	��I+4�t��=q�� ,}ɧ��O�A��e�}� �e�ጵ�W��]�k��y�Y?p�7W��R�+�3r�����!
�!`�`��N4|�r��<�6E���b
F���v:�+� b�
���Ɂ��a��r>f�
cJ-��Ʋxz�A|��ˊ�h#��'fИ�(�YY��Y�==Q����N_���0�	B�4�-�yoI�tTrؙ����㐖W�q߉�K���N�`�H�V1���\ķ8�`�����ǆ������NuU��+��x܏m������J�e�OT#��_\��cJQ)[��Fڬ}���3e`��o�2��P 	��;~Â��:�8��ak��.u�s��0�cA�tW�ԘHQG�(�"U$��_��%�B���<D�Uaxr-�nkU�>�I�S-H�z���GX�(
�Ak��<#�R,~�V�,h�3a��|�:�V��Y���kċ�L���kH1ת����+��0
oɳ�%=�V�;�&�Y��1�s�U7-�̪	Oy/���6?`�A�S�Ó���5�<��<c�TE%�}�	�W�7����9g��w?ci���9T�ڮìS{l�G�"D6v
�+X��ݓGk���'8��n�M�uV\xq���T�*Y��EL�N�Jc�����0'4��fČ��,�1j5�'�]yʭ'�UgS��;�y���^�S��_�/�1`>��	�}o]Y���v�	{�?c݇�^v�Β�>F��n�BA���yX��GF(K�C��6P�FQz���/��l���xgt��3�#�_�J�B�܅��(�U��e�S�>�9���V��6|Yxd��#T�e|ٴ�/Z�M�n��6���
��۔N����I��
�;��y+�Ls�`X`�޽���y�{�qs�O�p����5":��Ez �VK�'�V��Y��2
{B��me���.���_ ���E'�(83M�����S��n�;41�G%�)1��	���,F�h�^*�2��q˗��R�lm-='əF{m&�K���B(l�+5�S $H4qe��n��'Ed�'�OM0.���w]9�ߤ^�I4���MV���݄�l����R�'��B>�%ᕥv$,��i��9[8�4����嵴�q�b�ύ�Tҋ�.��#˕��$��#A��`��*D2W�V��Jc~���k8q�j�(�7�LQ�?ږN�U�i�`�y��g���m�������]#)��aux��Qc;��"��Kg�!״
`�jLI�;C����UQ��e`e�Ѫ�(���G�皧|�ՠ��ۺ�Sa^���x���'Z�9�w����M)9�3xs�G!��b'[�=�OT���dW�31;V���k��h����GK~p=��J~���f��Bߞ�&Uk�'�1�X��y�����v�H����?~p&���X;2ЊtN��]5=�wl%�[�g7��J}�q�28hG�=4��.��J�{�r�c��V�!�q�KS�xb�F��Kfi�z@ �I)��F��`���.�Lw�l~/����"�\�n��S^Gj��v@�w���k\��Ϝ�E�_���9�fz�w�@�4��O��QIb]�Yտ��k|76�3��\�``��R���A1l�wڽ�Y�
zA5nC ������)�iK9K=�<;���ȇ�� ��R�!Y��>��23�qf&N�R�f�VH��[*���E,R�tt��o�@'��՛�^vI��u3X[�%���ҩ�Ss���;�ծAZ��p4�0�,9I��
�Q��+�!Z	V8�Aj�����p�\�{������"~�jn��hr��T7)�R������U��J2�2.��j�K���̤Akǈ+�!8�EA���~/�e֜�?�0a� ʛ>�G��ͫo֐?�"���@�pLEFZ3�HK��)T&��n��C�||�j�i��TU�$���.�bQm�DR�4y�
��R�KHGK-s��h����W����-u<6���l�ͫ���O�W���|�EƲ�C��;f��	ۃ��t-�9���$�  Q�E���8UN��T����]�	�|�c߶ּvj����<'���@&��Qa��l�$c�����C��v	�Q�XjN����� #����G2���"��������P��Z�Vq҇7�af�C��8=��rgJ���� �sQ}tR�Р�i��Ag���Gƃx�eʅe���;�;�L=
 �߂��~=�@KY���l?��m��)z1Ѷ��4�F�:�wd됚���6��Ѹd��Qr�0�Z6woȑ�����f/�C�n��uD�N'7N�$���|�Gm�x�&��dK��^���IZ'�;~�'2�x;4��e?��-ɒf��(A7�I�H�m�gcx�7�����Ms���G�{7Zo |0@vҞ�ZO��M�ٙԙ	8Ղ�O��ିJ��Y��	�rp��&f+d-sK4�����QH�i#^'|����3l7V-7P�߬�$���'�ޮ���R*b,'sp�1ܵ��š'=#���� M��OUö:��3�&+��U����A�"�����2��=B�?<��!��P��Vo�0 ��T�}��� mj8�XG�<������@�������A5JT��[y0�ʗp�s*�� ���'��G�
�9�%�Z :�ѥe�[ڶҎ����{������,7@INa�ɩ�k0�F���A0���"y���Ŭ�)�p��SC2L�:u�؇�-k�|F���F����c�n�H�G�����*Χc$"�[��⨡I��A�x�+	�iHǁ�3Ŗց�;M7�,,��!�TGOe�*��yn7\��x�ӾM&V�sGD��)���Y��|�ڣ��`��X���j�l'+K(��gvC��g�s9�A��Q�����hv�����Ш�����&�łr3�39�0vV��VFЅ�Gq+d��g���|c�pv�EB�h��|O� �HQ�x�7���˟J<=^ۘk��t�N�<c���.��ahqrΥ2{7��V�hu�����Eo�1q87t�׫�I׊�Ս+���
l7��j���w���4|.��cCF����I*Y��X�oe��}���C�����?���B-1����A��� �^(�2�0�VM-�r�{m����rey�JÛ�(ଣ{�H�xQh{]���с=�f|
����w`Q,՞ZW9�cϒ7�팜�s����ݕO`�zuꬉc;��P�*x|lo4Q����qC�L��{������pW�@(�oI���}�ʄ��n�O�`�ksV�=B;%:Dh��?ԮM�k�l�XmG.'�Y�Mz� $�@A͍3��;�PUL�����-�_� �ٕ�p5�t0�ā�®�,�:O|Om`������F�����M��J��P��iLx��c����Ţ��S�j@� 8U��Ta�^37-�ͫ	�ƥ��E�	�)�^d3w�l����#�o�i#- ���1��2��4"��=�P��q崖2�e��ܹ��M�'�ȍu�(��[��\x�.!��-g�9"���r:��)a��k�9�K�)悵��	$���$,v�z�Y��=w@2��Yx ~S��]���2.]^K���v	�d�i����v��
Y�k���֔cg��`;5c�I/n%nEׅ�|�{ś{,37��wGn���#�~����`Eܔntp�9TI6����IS�aؕ\�=i�r����Һ@��@��O]�����N�q(J�~��q,�Sg�E�w�;��kx�=�G�?���8E~�B�ŏ^����0�@����
o��A�DɘC�d����;�*���(խ�̡ys�IEqL�2M��\�C���^1֖o��jb�І�dP:@�`�k�HqX���ݳ>"�l���9vڎ�(� �y��.T���v�����|��$QB+W}�Qe�ϗr�;��f���� t>�
h�a�V|�̆�T��DvH�Q�Eյfr���Q!xx���јw-ܞ��|
�p���U\��s
tk����\)\����۹��J`:�T��Ҍ�x&��=W�i�c������0��M/E}8ƫ>�?m|r�c��I��j]�"ׅ_O��"{eV�	��P<��T�Y%&�G݌�3�+-
!JF�P�I��}�,u�M�df�;���w�D��zп"'�(R��"F��uF��5�K�y܅?�-i�|hՔ�0��W��(
F.j�`)@� n,{�xF��u[
�v��{����w�>��5m�!<@ x���3�Q��*N�4=�fڃ��s�he6��cҞ�t�h��!ٍ�ƹ���Z"����6� ��4d�i9ڡ^S���_�эC*�h��b@
Va�Jx3z�xR(��BP���8��H��ys{�{�~�=G����,�'b�_ʑ7	r�f e��XŦ6%l�4{2�p���Iq��M��$�۩�����YjT�|/�cߦ}��6<��>��ᐇ��F��@��
�*h[JR��7S�W\�
ɑ���h�s\L*���
b�d��27����n�-���L��_�,{D�U(��&ߠ0�t�>v��D��p�}��Xj�)>�t8|H�A�Q�К{ya ��xnyJ:嶄�����؄�sz��!RI޺�:SڋG�:�e���ָ'�6�*�z.n݋>[1��bp?%��9߸��zX68\o��r�6�$7G�0��UԀ�d��`�ß��^� ��+|i���K�?��99���ЊO$(��:�{��b��o瑸�V�c�!�5%�K{{f���g �p� kzַ�������c���#%�'$�	0��Q�;�2�
���ˁ4�{�
y����!븣cᯄ�uEi����]7=[�[F�İĹ0���3a�L��Rm&�T�����{�ڄ.�y�i�[�Ղ��f��w[�;�
��ۉ�rA��5���a��n%��|=�kh��z�b���J�{��%���ʚL{j��k�u����h��x`L�U�"RϺ)����u<�Q��0 ؆9�CR��yH,1QI��s�/#�38�y	��a�|�(wܻ�d	��s�꭭�*F�h��,J�Z�qÉ�	6�C/��>h?��e���������"�q���c~��4���[��䪒!4�\߮�2+�v.�|_9ȅ�Z��"�Ȍ(��Ⱦ�[(�p"n��5�d�m��#�=�\��=�>Q6��8,�|��ZkFP6<|p�P�Xwȯ-��2U�;��p]6�x��	��8�s�U�JM E>��5�;��9'*I�cvi�����\h��M! �AG�2�~���B溤��>	�),}Ĥ�^ؐ	����h�������)G��t���>�ܦ�`0�W(V*���\	c�~���Qó�*��������%)C�\��-��r{�8@�ů	���Au�wz"�4�s��l8�>N\4gi���ɷ��%hb�т[��;x��w_I���KF��b�Z:5|�����O4��e=��MŤ5��3�m,ۂ�3�^������zN7#�l������+��.K�;��~y�%�ޮ]˽5�� C��6K�La=|�V�ӭW�3�"yA�>�%����<���3k]�2��������ؿ�]�OB�;Y�Q!�=<����x?�c��X<Bs�%��|>�ޒ��dÅe2:���b��Ry��$�bF�K�}rx�)�s/l��G�oԞ =�V��� ���]�5����O����;N��YS�.�4<9-�.g֬���͞�̊��Y֣.+�=3�����t?����c�jݼ��9�ߝd�<�B��U	;"��� ���Qȓ�`���*��z��ՙK�V=B��Zh�ռ�#�W �U�Ђ2`�q��TP5�z��#��WF_�nPY�m��'aJG��0�g�S��V�'MB�C������펢!��1D����>Y�P��W�O�G��d�O'�7ow�'��i_����E58l_K�~�Sδ�W���KmyQD���4%>5mB�m��Z݊�Ub*؏e\���x��@��qğ�<�=��N�9R>����Ka���}Î�#g�,{�������h���w�B��̟��rfIb:� y�۴��9�uT�U��T�zv[�*���
f1�3&rW�*m3�?�I����kv���0�o�	Z�~��s�s>�0�4�(Y���1f)eq������Q�_��qbtr�5�6e�0�s��<ゥ�Oֈ�S������8Cb���@	�1�X�b�Z���Wޡ�a��_oC�#�߸��̙5��ĸ�U�3�Y9��]���ݭ��G�Q������n~x�D�Cdf=ƣ�_��,�HjC�.,��!���^ ���o�WZN+��䅳��mjվ~�>�XV�;�������y�ȓ2p��F{.fK�ψ����G{��t��%6�L���'��A�of�%c�6 L����P�;6f�j��ͶMx��F2顱ԕhTE�՜L6Qh���3��ս���Nhi��ǬN�Vk�hl��$��5�_��܀�<K˒��_p��E$APA�a�'��ϊ�A�A�M��
ϣ��������;�|���C�-R�V+�k���~�=:-hX��⍸Э���{y��Ƅ�c��(��것�^����3h�x9��7��Uq��E�gu��f�!�.Kg�:>���YJ�D�^'u��8�� B�u�B�*�,��\f>��蘆l���V�3�Oh��7R�����H�&D��p�ƉJ�>�l�aCy�8�_^��M
��������Ҳ��r��(�?j���M���`���$�)wc�S��b�
��*�p�7?(o�O8��^
J�XT�U�&��?����s�lne	�!�w?GR�\r!�{~���͇,�M�6Ri�-W[K�� @�3�*�"yVm����6�2*?Sg:��Z&��3M�/�2h��B���Fݢ��h�|�'m������;�3#x�O=��h�|��V������7����7�`���~AK-�h/Ƙ^Cn���O�_4B������3�M'��V+�_z-)�lu���Y�E��- �*6Q�!�K]w���(���틜>�wK�J�`�4�G;ɣ���m�<'�| ����|1�ij|����-�I���Ok��&�oL�;Q�
w�7B0� 4>�p��;ɚ�{,H��V��^�ϔ,2���$��	N��܏�X5aL4y�%�C[�R{ۿBU��=�"����v�6}�-�?.>_��ɞ���$�P������K���[:a���ԅ0IA�.�Z7���m��s��'��W�E(�m?�X]UU���[�:2w2&;�ǅ�W���abu���\Su��lL��"��T�:�K�Í�p����.�$�܏UM��V����l �'�Z�֋{+�3b��p�L)ɫ��Cu?h��f�2l	[��gp��iD��>O���@w
����YE]�F���h)�f1KK�j���u)�
K�#��^"��+.��3]3*�`�\��(ܟP�XD�&��Pk;Xkq��4�|Wk}��N��˸��sdoAj������Ъ�?�w�o�����j��������e�t �٬WJ݄ �͘��k��Za"!�5�Hu#��GE�3]�k������.x�v�ͬi�GrbE_�߫�����s �xoMC厲�2E%� �~ؼ��Uq�W<���a&��w�H���^�6]��?x�~� ��d���+�(��M.>p
A�� 4K�9l��:3g�9�����/���L9d�<K8�ۙ�,�u��o�2�������,�f��y�B����+��m�[��Ejh��^��:%�;�(������V4VcVm6�X��ߓ�L[��E𑰨En�+WI�%��SA�qM�lBqH��`�['��'M!�xF&T�/g8	�p�o�^�J� |%=�70(�Ϳ�t@�넲1���%��(�c������ͱʄ4��6YV�S�߫��+}���GA�y0H���4�H=�r�H��d�p�^š��2X&Th�C��љ� Ӭ�4%xO�w��D�*v���F����vh2���8ڮ؎b	�)6ҬKl-��fK���H�H�4m�E��.�߼4��|��ҩl�ӗ�
��0� Y��'/5������j���.�� �Z��!�%i �����	�og�f�n9M���gեZ۰@D�>lSh����x�U�� ��	O߳��}'���D&���kE��j�`G�����jȜt	�yՊ	��G�A��+���6�i�}��{b&�&��(	��w��q�,gҞ/��cMo�<.��qE�Hh����4�����}@���y ��`fU���'��A�3;�΢�n�@
JoƂ�e������yy2Yxw5��
r�l]��'Fq�0�[0�f��b�������]c�(㉷�:��$lծtW�S0*�7�S���;��fO����<T�Yơ�V��׆*��C�)z�ʕ�`ɹ�Æ-�1�K)��׮U�A�,�M�ή�ޘF7?���S	�6ٔo<�ޓ�ͱ$SpƔ)��XG̓�V���,�9���pj���r�y�~�1�)�� ί��,s_V��������6��U��Q�H;Ӫ�5��$]�i���I1�����7�xe�LdCD+\$�|ɛ4��k�6뽸���z���݇���5>��ۗ�X&>�M����U���!R����1��G���)b4�)�K��� ��(v7k����Dя��oE�D��]�\V�g��i���x��ͻk�PJֵ��e�0�U��T����^Cog9�EM���?bz񎒒?8�ڿ+?">�U�I�:���tjت�э��?ʻ$�����yH��縮�ufH�����	)��������Y=��hn��BGӤ�Ud�!v<��a��1�&"l�Z��"^+�5�l��&����Ko�x�%�J�D�ƃ:ª�����kГ�L�t֩;�ϧۃk�`8<��	���+v�M��S������}�Q���(f{K��%��iQsS 0bzIh���*w;k,�1��<�/�Y�ZY��t���&'�;����"/���PS�F�;�j���v�r�����O�v�]O�i�lUٞ��/8���Y��^7Q��"�G��F���t��w�,�,p��H�5AA�ʡ���[��^4�w/^f��ۈ���2ꉜ��{1PI�!ߐ\�WR�p����0����u�s$���z-��i{fK����W���!��'�Ӝ�M�P{��p|�A��s��IW����?u�^�g��ܺ؅�^Ư�<�mn�U�`�!�*�{"0���k��ކ�xT��!��n^D'��mM��H�t����g��W:��ɫ!y��zc� �V.7��u���_J�X�nͷ��D��1�qh�^
@�ҫ�`�׍fCe��]�a��Ќf���:`��b��=���������ho2D	���FI��륾9�� ʲ1=D�฻��Q��n�M�Y+h�S�e�]o�C���;ܿ�����)jBw";p�w*�Wk�,�A�׸˰��D*�s����mg~}�C�]�a����ewH�K�#�ު��|�gSJ��UW0���u7��v�������ݙf��͍�B�����o�cv�U4�i��YRd�D6y7�X��d$~[X����	����	�T�S�d#�J�})�X`<��$����=ծ�9�]K��SN0J�����c��R�iӆ�%�)C�bN7�㣩�\�e,	�d�#d�/�'#��?�X�����+��%0�G &؊��Z����M8�G��&�!�0W�g��_�T�����3l~H]}��X�ѷ���,$�.�;��CÙIⲚɣ�h��a��F̅��n�pj~��`����G���uLG�M�hYgS���1�Tr�u㎣]ߙx0h�2\V5D,;�����4����F�ݺ�WG���ie�d��:���M��2E��>�0~w�\ݤt*D7��΁S�1�L�>\�z��Q��E��T��A�L��z����҄��a���9UM�����ך�F@�U^�?���X!_$���u[�b��:K�<Z������z�����֨~������7w�Zr##dHiɓ���/HRɏ�r��=���Y��8O\���%��u�Q��Kw��anN�#F�YR����8cgx��J����We�=J��ń����]c�p����@����9���e�nq^����\�[��M{#b%�z(��!+ɛ��a0�H޴��݂�别�X-Ut��T3Jbyo��p`!=�e��c�CO?���̀��C̰Ȯ�`|���L���������f_v|n�@�D�k�
Z�@��st;��h�x]���ҠJ<r�.��g;y��)���TgH�U�)�e��7��9��e;_�W0���q
��~r�x��/�7h3LO6���@��;: ��e9��+Jed)���(��1 ��е�>V���[4�0(�S2���hדl@�������!�I�Hش��J�͡\p���������c��7�D����=�:�I��89�O����@>���V@5�`��}�]Õ���� J7����N���]j�y�9,Sa��nX��̫�ܢElZ��4PbFG�
��͆�T��F/뮉7*3.#8����~o�݉5���#\s��W��w`��^��9�B�@��_F��ܚ<}l}�&�TR�3۩��l�z 4F<Ak/{i}$I��SgO�i#�@6]�֧��l�~<�[&���$�&���t2�����:���	��'�`|)@�1e1��)�1?B�G��p�Q �S;�8�`L5�0�q�9�)�A3u����	訡�E�k������H���-�4-�[$�H���^:f��*F�ڜ#��v�����MVDN�K3%5���!+0���Z�I�:�ofDbq8�v'�&�ʬ�|]k`�N��Ĉ ����n֫A���������zf?#)xq{2�e�*����c��f��˝n�����
f�1���p�$FS��/'+[y�I�
z���)M�nV$����±6aJ? N�x��Q1����x��d���s.�GY�^���;Ti��rgܽ�9�t�K�i^�I��������^Ҥ�'���\mT!nL�k�j��9�i�Dl���g��>M���:�"���X��&n-��kӛ�x��rj�?]�!:9��j��9L+^X�xN^u�L5�̲x4��?�pC���O����@�&�Ͱ!ȨC��?���D�{j���!f`��Nf\5&k����AR�5�������BT��kȻh����n-�r	��+ϕ�tR5�dT�2�;�h�c&t���5]�8��R3���~b�D���"N����Qh�\���D��,as �3�7����8���)�����}��q��p)����AlA_ubg��pЖ9h �5�����'�=��T}�׮Ϳ�����a`����Gϓ1'J��]���]��VbM<��;�aS0&��Q'ݨ�V����9�df�d�^B���'7B��v XD�'/Ԇ+��>���
���)�4�(��_߭ �Do��B��]M\p�����q]�gq O�i5;������.r*���̄̿�^��a���p�H��$?"L�~A�F'��8,?���
�#��T#�i� ��-F�jֹH⪱�B���U����N�>�����XF�g�?�\�i�B�@� �@L���ҽ}<U�XS(���*ͅ����@��J[�����v�U��ot�݉� n����x��*���f-͌��@\`q[��(V#?��s��a���h���(�ԧ����j��M���o���Y� 1�=��
B�9^��E�YPW8���T�v	��(��E�'<W¹�ũ)<�.��J�IN�V��_f	*� :�Ӭ�.є�����+ckΠt� �VPBg�� ݆@�qF�TSm��:G��Be���,^B� H_�^�Yiل,Z{\��4��i&o�=��Ͳ٣'"dR� g��|J�QRX |��Q��c�g��_��v �����"U9�H�?0���6��n��>��c�����䩝�� 2{"���&��,�Y
��BV��O���z?�-�z0�k��v�����? &�]�)���1�ϗX�ԯ�S�2��k�ǣ�Z�CN��mD��ϊ�ץ��ݛ(��½�.���C�]�7�e�L��-�s�2UyJ��e
8^��C�Y��}������W^��o?*�����Ne���ݗeD��^�Tt�X3�$���&�<q� 4���	*�y��O����(��|���1lR*�J+���W�#9ikv������@���O�rT��O�}��
0�����0����ڐ��Z�U��i��ց>��h��
[Q��"9��(-	��O�ي>�9�r����o�"�vY����S��2Ҋ�c�q4Θ��Fs��B��D-�����@��B�+�jPWNx�fU7t���)yP��%!�	v+_��㩀�1�ܮ���M_ �>Z���宮"V�!2Uە|�J���5к�gF�aw�z�=	]�����F{���Bأ��$aS�~��f)��^��9#�q�m�f�1�����O-
(*�Nvꤠ�-�pp�0�<���N�Mr%����]O�QI5���,@�r���$�K�8.ʜ��ϴ����*�<�P-F)�I�T.I��A�9INA���S��R;3a�
���] 1��&�tE�w���Eys���c���Y�Ekog���,rU�L�m��q� '�5F%�_�z��Ni�֙KwY����)�N���9�P��bo� 2�{�� ���T;ݿx�˺ۀ�6+kѹL��KΜf�C��R���F`C�9D�y�,���:{�Ϋ1�Z�HH��7�`P�o[Y\=��*��Xt$�	ެ��(2�=����]fPB)�.�8u9u*��x����-�ů"sh�H1	��p�٭ |yӒ���d�ZME�t�|ݣ3��E�/��%)EuP,qν7���H&��Iţ� �IUN�'%�H`|�!���ǂ���Z��Q{���������&>�V��-	2����5��A9@�w��s`vdAu<��p\�;A��"���/��F)�y}L"�F�`m�ͮv;����Ӑ�;'�􇹩�0���6�F�(��tCJH�{�d l^��h�ޫ��_����4�nC�R��xfa����q���v�����0��@]���K���1�~����B�^,4��(Q\e=�67����C��;�L�62�a�m�KH�����[d�.��
H��%RTO�fw������F ����~��H/�Rj�麊�%�oP	��������6v���R�=j$���
4i�t�-�R�D- x���/0���F=kA{/k�����
	 ���g���wr��EŬ�W8�4eOb**E*8��
-��,;p���O2�?r?a)�JjiC�qN�_�6�NP^V*�����r���e���'g-�;s��8���خ��[$U�!q�?��.�H'��h��i0~����+L�"�]��C):�I_p�f�&	�p#Jzʢ�{F@%p�p��[�hL�1Ρ�&�-�N{�D�ҀPj���c rD`�e�LܱA�bËN��(���l��D&M��0�k/�{��*"��}��e�g��l<\�Ymn��>��Ϣ=Ȍ�@m�ˏ�"�cE���1��K���^ɦԪ}��G ��6lr�/3SW7�z nq�ْ�u_ݕ*����/\�~�އ�L��+W~b�Grc!�j.,�/���������Q��R�n�i[hjxr��[ۃ�2jY:)�<�x����QRD�U^��eǂD��6 2b�ĺ��*dU@ޙ�_kC,� ����] �����	��bH��T/�a�//����}�ٜ\`jۤe�`8�X�Ud.�$
��9����_��<Bl1��mm�٣c�fh�GPp1��!�o�Tg���_rѐ��*xZ����%i�f%ĵǿXD]�2,�f������u��RK���>��"*��eT��+�~��c��v����� &�ʦ�G��2�a'*��ؕrAƨ�;�&ZD��Y�
kL��l��2�V��"hS�O\���0�_k}V�@:+���i?4c�%���.L��7u��d���f�DB��!AM��ioV��W>���ʗ-'L����n����JC}�� ��㟰K_k��E\��u'ģ���@�
I����^�ߕ��iR4T}%�����xN���З���=c��ޚ��{ġ�]M��8�d���z*��(�$�Z0(�a���;����#oc9�w� #�¥�6h4��;U���ɹ�0�>jv�ÅK�l� ���gv݂�e��U`�h��L�	�7�犖j����N����n���L�Mh�B���^W���vUP�l�λ��p�#<I筙'g�@��49���MRvjJu(-]�p��M�����JR��]C�^4w�[J�7�p��erQU-��C�1}3yB�>�y�8�!�Î��8�����_5%�zq�L-_������, �J5��H�ƈ8�;����(8�ؽy���@ �א���m3m�]�o�j76ʾ�đ����-�$��#���4�C�Es�@���*�{���<�ux��I�١��Zΰ4�c��b�ӛ4�(W�`�K�č'^�Νtl����~k�n��YR
���D����Z ��h q�E��vƦ�n<��B0!�T����uItI���ː�vaZ.�T���ަ�Y��s+���p�t�����n�BR �&/fcGy�������M�ʺ|b��z� Ӧ�e�
�
��0!X�>Fa���#6�O��wn�>�����N�_�&Y3��o=��Ğ�6�{��|}�01�.6Bx�IzeN�>�����!:��vL�5itW�/;@��[D�P�Y�[��`��/`��b���+���z�u�Dgln�C�G�R���k�K:'r��'���6�!����:����e=k�6,�ը�mVR�fFd����w�["�H��/����:�x����f�����_}���I��.L�\S��)l��4���Ӟ`�sUls9zY���;������@=����5�R\>Fo55��/D0��rn�5����|�`7���GQ8�r�Y)�f4}��!�0����]
����$�$�s�0!�c�rd8����~l�u���G��Uˇܹ��8aHF͛}}O�5^ϐ���?�X���I�g�7I9��c�γ�u�)+,ui\+�_������!xw#�D�jqo����I;{~�#@�[�&e���<�WZ?A�fP9Z�`�oq�$\]� ~>��q{c2�&�僚�5A�4/9����I�@� �b�d���+��������6b��E�(�fa9?���["�ф3���4�.��Դƌ���w ��77��������NwNZ�	�y�_ToA�~�3ÐR<9s�
�#mB^�����N�t�����6!5��M�~i8�����NoM��4a]S2�$�¯�����Ή��.]Z��H�T����ߊ�X�<�1K�H���YF�e����nZ�l1e�M�ck>�P�ؽy�����:h¾b��>�b�=7��_��6�n>G�y�L7���5��j���옔����S[b[��k��_�;��n<%���[�Z��gKE�k[�1���%�e��/ޤ��fM^��Ev��~�f;P�jҩѻy9V9��e���$��壥'���¥)�k�T���"a��S=�$i`�aH
y:��������=�5&-Y�ܽ]<��$�l �A�Ï��}�H��]�������C�6�V&6��׍?ȅf�,/C������P������u/B�N<�APm.��J/I�b�m2%�ӫ��=�6�Ǿ��(ٔR�#������� 9��n�KJ��:��!�T�Wвn�D��H}��?�Hm�O���!<��>���<?���5��.k�6\om�^ޠdE��(��D+M����	8P�{R���8^�1J�c�<�[�@�&����x׫�&y�	.9�G[���M:��}��ЮT��F8O�<�\�na��G��llݟ\����%�v��ȳ�u�Jƒ�/I&�s\��}�;�w8��[��r��+�v˄�z�>���t�K�k��ܯ�b�T��w���V!�3�z3��]�Bؐ��%�ߎ�������  �Y�r���i!�]ӵ�o�9�6tZf���J�	vV���w{]=g�EN�!v� ��d�G�qP}j��'?)���X��C������ۑ5��sP�~i����ctY3'R�L�=8�M �Ź�2t�:)pz�����c�/f:��X�Lu�~�j���#cB��ô?ɳ��g�s��e(��?#4�U}���@��gz�n
���G��0�4Δ�AJR���Py��� ��R��U���G���'2�N��5�Wz�\��X|ʮ����J���6XDx:b��a�H�J$��V� T��/��M``�f��ZKT�r��X{j<�=M�;`����1�4����{���0p"2�f�N3�Od#7�L�}2�5��:%�6������<\F@ )�9�ub�
�Ոl���HiԿ� �b嫯�s3�w��U�p��e�k䭝�'��&��?�h�5�Ԥ�T�\�7x��)���R�o���iͳ�2��9&U�|���w7w����쎈Hג<��?���������6?�� b[\!i��1*������ˀg!8�ACQX*���)�8�X����|��T��O��9�}? >m��gl�����X������x���.p���9�����G�k�6�	�T6��8�+�i�~���h���2T^�w���P|f�"93ⳢptWF	���R>�%NsO��>�l���>Y����3�f6���%�c!�?�}h��;dii����j�Î��BN����D��k���`Z<wx���t�T�8=\���K���`xU�Ql��;Kt����o�8���ou^|�������z<�?0�'u���w�>o�v�&���oj^�ΆGmאx�0J���<Ż��[J�{��T�E�	!�_��������9.7S<vY1{��6&��]�k�<�O�̒��#�b�Ԟ�M��n�)���!��Q��y�Y�w�-vC}H��u�g�H�#j'��Uo�>J��5�e\�el����}��;�	q���c	��(	�,B��P7�>eꝼ�Q�鰋�GP��EoHK�J$��D�6���37>8.�߬w\��\�妍)y4^�[3Z! 7"fDE�g��`timC �(����2�yK�v���!���� $"������֝�(;@���+�/Y��.��x�*��@�r�3 P��m��m��<�ZÓ�:�.��s�&�}���`S�Ӌm�����RArE�4���d�l�2��$KO�R��݌�/1Z*]������Rr���k�33nI�� �i��,���R_�'Q^�bD䪈�[��O�#�!&�2��T\Q6����KT �r1�d:[0o�B��Vci�.\B�7�*B��O�XȾEyaw��A �!��9~Qp!�m�(��%�j ��LZ�V�U�T��lC��g���.oz!���c�lr�w=6r��L�S�M��l����!�(W�L�!V��+�T�<��Gb�	�����*�AI��l���zT��0�!� /2�ṵ��_}
���Y3hD�iXǑ��g� ��4Ȏ��U�Hn���s6��d\��U䷓c�ŕd��H�G����@y��|0�{�NӇ�������w��Q=��Cⰲd�f״��@=�u<M�N|�Y�q��v�
v�q��X��ؽr���5���q�r���$7��F�.�Z���ʩ拔"H�-�j�V�P�$�e�[���r�0�+���6_��(�Ig�@��T��) + �%k���|jT}���Ƒ8���Y��D� ���&��phu�3F�UW�U���v�����\�M��I 0n;U(����C�i��q�k9Y��´I�%�W���(�6K�H�8��g#� ���o.�J�A>�����d���-(8��Gzu��>��'R��O�M~��P;
tL��V�M��H9�$�db	R���·�/�l�F<s���c��lLfl�ta޿��.<�ҢD�3ˣ�^T����M>���y�(Hi���S:��`eKCu7��5g_p;�*o���o�+F e�{�+���_���x�%0�S�y�@@�r�՝��u ���*�?��
���^��_�]�8����Eu|@-���D�2�![uh6"�s֊#����E�9�2$�p!B�K>��₞�c0�Z�Q�$/��rq)2�؇�A?_g��~3~u����G�i`����BK� ֈi�n�*�{�O#e��`v�ø]jQh��<R��Ӻ;.�m6C:sS��i�r��a���lJLZ�c�x$LM�-E���Q��Ŀc03I�֟;�W}J��d1Ԭ'��
�k"\<�RB���瑝�� wh�o��$�vg��l��f�zVt��
:�o�������b� b�\s[�C
��E�զ8h���X����4�@ì�[2.V֍L?i�%�?E__��̐9��<j-�p���A�0րA�'�ǈ����t� p�8֠_����7�vr1�Z�x��nj��O'������!��r2D=��O�Be��ј����`���O�C��F���`��d�e��*ִmT�� �/&'�nn�W���1=�Уv ���u�g�6��C���U�����aQ�����3=�as�X�������p�J�ސ7������@|5Gڊ|������]j)13̙�n�|��rr�.
]�x6>�GĿ��0�57���9�ʎ��9Ac�ז^bf/a9��O��.(�'�P4E�	-˥% �<,���l�t�����+'J�e�hn�h��*�AP�S�h�;<��؏��&��x�L�f>]��)9Y��*�1�a��KCh{�Os��tM��b̔=�V�8Z��f�'�
���[��8G�W�Y�T�T3���Br��c�ĎYQ���;J���c;�1f����K�su�Ŕ�t����y�T����Q�N��۔��Y��s?k�����3��f�AIx���/������J��x�_'��kJuZ�}��5+I����	����r������Z� kIٞPh�^��K3֥U�����e?&ۇ��������\���~V���ڎ��!�gl����z����HM.�
�E�:��e�\X�8O�.��d�g��V�]%�FC��̒$��� ��E����7�=Bk}��w��5j�w�6Ԗ>�s���v[ޯL��r6��n�h@�+�Vǅ�Pk����k�Qڔ���*�m$H���	����[�[�(�W�G3�*}�nNs ��ĉ3�Ri��_0M$Ќ�D��?����ؑ[���Ǭ'��7B�U=����$~gQJD���NMa�x�y�N�-��R}+���L���
z+w������sM_C@�5w��y�Π��b�Î��Aw\���?͗R:Ԕ��m�mt��4�/ܬ�U�s_�`�-�+.΅:��V7�Kã�@Ʌ�w�j��[���%N�N���F��ݽ�:���9�g8D�X�.�}	���\ �����p�F\�D�d�*EMF̆�����J�i�UJi�8�B���w��RgO�a��o��8X�-�+Ѯ_b��89��;g�c�}eb�Z��Ǉ��2��9��_�gCd<��_w�E˾6p�y�ߛ&64Hu	�V�:��f��@�ר0r�'N��ˡPe��hHƧz���ɑ���e�<���:½O��xu����	�Gի���1-J9H� ���x��A�ӵ"5�L��}0��i8%0�Ǎ����o6�'��~n��9��D�ju�#��:y���_�[H�(�g'r�x)?zM�np&8ż���^,Q���23�o�:l�.]�bL]����5�$#Nӡ��TB���P�뚬���p��{�$O��9�2m�jU_�X�t7����GM�#�"�;/��j����XzSo�|~%Э����;��Jj�bUC9H�ܪ�K���:������pɥ��%j-���©->�'�1��#�%_��#>����`"y��74�Cf��V+ݛQ����C��<@trY�aqb&����Ќ��*}��I{C��%��?B� ے���9msj�'E�Fe���8Q��2l��ܪ��;C�0������%�T�3
�hZ-
@���9sݲ�KI˒�'���ޑi���,��� J�~���4,�(*e�����F�
N�I�Ia�9�Xۏ����?�dW��Պ��˗S�*2XÙ���.��1�izL�]Q�v� �AE��?���Dm�Q�q�g$������˝(IgG'������ռ�@��1�X���H�N�{f�\n��"K;lO���B:�� ^m����M@z?�K�%��{��x�h�V@��9���Z̖%X���ퟒO�OG�b�9k�a��~�p��w�|2�lB:U�t�?Ɨ��[���L��І�S�`������Mc��e��s��Lx�v�l[��lh8�]+RC��٬��-G����&��J ��ѣ�)B�+�w-,|y�H+�ͷ��uK��>��~D>}6�]���w������U�t}�>*���ʝ�M��G��6��!D�B�P�:��g��_�U�0-=���2m��R��|1��M��*<R���:2��Ur�޺H
����D��>`H�݊���Z!}ݒ*��St�}�V�Ät�f��϶�}E
+�m�Q���n����t-';X�Rϑb*"Zz�|��ªi٧lך�;��z5�,�碖�1R`�r��p�m��a�撋���E��@|0��oY�lznh�g������bs�����fb�0�t;��X�m��
T��):B7pDgx�O	���ع�7�BS�A��y�_Nj���N�Z�1`Əh�;^���Q�`Vނ1�3�ؼ)�Ǐ�?��a&<l����"�J�"��V�q�	vhc�+���U���sH�&��V��ns¶�[�Y���JN)�kVdI'�(J/���9Z�?&�͞��o$Rs�Ht"�r��-O�o �3�NN��;ݨRM���G�QD��M�\]yM
�K���Go�j��jB>$�::C77a��.A�d�vٹ���xɲ�a��q�� q��rhH�?n��"?Ü�0�5)q�Dg�V'S��!�����ۆ�+{�[��Y�֦��6)�o���a�����U�m��R`h��ɨ%a������� +#�*j�W��9T��sN%�:����@�SUt�0���+rv�҂�xɎc1�����zR��c��%0n���L��
o�	�כ��{��Y�ht*C6A�+���;�h~����kP"�2$��o���~It�h�:oKmX��%��뗿�X�G@�?o���x��~�����ȱԜ���e��S�!m�NV�	�~������J>��+���ҳ�F��H�1���\6E������~D�vo�L #�}�!�Wj�xS<{�n��vr�����ؔ�-�J!%K�Jl��d?�h�wF���ؒ�A(��ڈ�
�]a�B�����U�H��-���������^g�ZX.�V����AjA+Q�T�pb��KvӜ����O���FzV:��_J%I[t47�H͐B��F� �K�4]{gCP����t1x, ��<c�&C=��±z��
��ó�J�0q�������2imcRF���w��n`$I%��ƚ*� $�)���۷�ZΙMV���-��S� \�C��d�M��]�.�=̵X!&\,�"��?Q������eJ5���0M���PV�C�YKh�e
/�#'�'T�JL����&0�T�2���Ko2?z��u�R�7��YFQ����-T�T| �9I-Y9!u0-n�m�	8�/Q*��6��:�9r��H�W+Mᥭ�g��9� �����Ɯ�Ab/f�S�%$_�j�[�?�h����d�([�$ �І]V�;�R!�|a�;/���/F�-�Q���.�����c��$���L��/�VR=e緰 �^��M��!��İ�%`2��W{mM�״�b�>��Â��n?��u��K��O��:QBѻ);�������N�����5!��S
�kD�X�^�Ғ�D�D}� �.�-��#�h�|rFFy?ܕc�*,GC�c9�
6>pm�Io��:�n���A�G�4*�DB+��	4��Z��lhݬY��v�?gz(Dm���J!j��Σ<j�:��������h��p�m��:ubD#U��&G�0MupO1��t��>�'�z��v�$���~x�BQ Ǒ�*�H�A��q����c7�J ��Ǯ��ܲ^[i��28b�r��"��]��иVMO���6�A�!�o�� ׆->b�uvꢪU��@x�@�Px~(�����^�<XW9��&�fɠ�#��քEz��n�̔X[C��sR��1>�s|8����.���%�,������ǀ?��<Iʲ�����B+U�^�d�)��� f\��~;m֓;N6n;���*��q��b���:kl\bP��A{4U=�ዏ~V]�+�"c�Q�U�����;�J������������t����f���Ѳ��|
ջy���Fz�5�8o��E-p/�9�2�|�ː�M��[��F��^kSh�d@9ݟB�n��L��u��WNfL��B����N��4�r��o���9��?�U��k�H�
xF$J���������N�7�F���3~֊8��s!�JRջ���{;s���fwJ����]�i�B9nS�$6���$o�zn�ŋR�U<��) ��T��+�8�ؒV1!d�޵��yZ?�(�({�V��K�6D������C3c±.��V\�ŕ0_�S�p�� c��6�r��$г���!<N�䨃�q��nm%�9�1���H)�0��_�[�M�Sɧ4׹��%+�ǺIbc�"b�Ջ:�Ʈ�f�����//����Q�
|1Y�����X�F�9i�*�`&��S>fM�9�d�t�f4v)�i+l��a�Rs��P��#J*5e=v��&SAY|�B��.�uhH�o�A|��y'D^��]�-b��juW��K��w� �E�����Y0~�r ��V��9��sh$C���(d���۔��Go�PI96��ρ�"��I~-1�����L丿e)#�:~+.������x��m�H����#�5*�p�B<���;�Ed"�<<��3�MD*�|Į��x]��!�*L.�Fۦ��g�3	�=}�ſ�3Ԛ	R�0�,����aC
�.������>�e�2�g�'Gk��Ն#�G*O����o*օ�i'���&�Im0GSA�~3?Zu<��e9
OP��ǀ9��Ͽ�	l�#��M���Hbx/i�8'sB�~�J�N ���q�r�.�!c�#������~�����@a���%\L�N3�7���ލ?�Sƒ8�T�s%t�ߞ�!k����?�Hn�E���yK��p[J�B����xL��a9��h,�g���i�*���/��Sd�]�קq ��$������~�gt���JK�UOf�"4��ڐ�k�<.Dಶ�9���h�Ȥ^x`�b�m���E�v�m!k�&7��Wh�y��+�DP��XB��ŕ/yYuB����Fِ��5dw�X�F�Qw��!��돠�M:���f8J�4��xK�ȜG�V�������z��H�.N�M�e�u?P_�����S �?���N2�2g1=yTG2m�,vB��p����ß��Ik���o
�A^��?�0�Σ���<��@+��al(�[�a��+���97�,�Lh�hx}�$%]�^Y���{�w����tL��VZ�	V2�M���e�R7Vi���p�t�\ό�+-s��<�gS�&ϴ�?����1���q�ks�LK`-��/:4"�˖>q���*�7���^�Vˀ��jv��<J�I6~����-G�6��F�=�J��ы�Nͤ <Ĩ�Ȅ�+�|!z=c�kg�AW��J���	ͅӪ��E���p��3d���wF|c>��9P�j��q�,�C�.�ݙ�q�|�g9��t�����=_�@y��wǢAL ��'�=�S��Ve����/-n�,�z8���U��g7��!Z�$z�pR�@xx�7��쐐�X��B�XbLl����V��5�00�P{q�@���#s�������1+ � �6�[-^�%�!����`��B5��n�9(DXi̜= "�7n��*l�x�7��Έ�rf������Y<�E��%a��1���_�Sd��C��,�z>��,`P&t?�����6���D��\}y�@���E����=wut�ɰ��1�̹��� ��$
�ڍ]��;c�>)�Ȃ�S�~o�'���P�x%x/��%�	~��������O0Z�`��cr��/����y;�N�xcH�ژ�D��/�v�[��w2�9�����g��$�\����:.6̯�W�{��n̴��a�O'ڈˮB��qe�,��F��ǒ{���X�*�~��1�>��9Ho[6.Zg�Ɏ�Ǉ	m��viG��t�ڎe+� ���v!�(�e��=<��5R�Ф�o���Q>� �r�u�b	��E��Q���s�3s/����O����J�p������4��.Ovf�+v��.����}΃����� ���4k�I�����p���[�3���,�����?m�P\�d������r��8,������B|w�N�#yf'w�1%SŢ�X��<�|�uDZ��͡b���^�Uɦ+�Xu�����	��_�B���T�P�N%�1TߕT)v ��+��"��0[Ϸ�Ɔф�t
m���y� �����[+�i����\��o���*"S��R�B\�!p� �+V��n�Y����v�G�R�0��]z9����C�T�i�^I�@�h|�<|es8�W�#j�����q�kOi�[��-���9t�M���~���a�O�X��^h�n8s�.NB ���(����J䠩2�<�.k�ݤ��y�X�Թo��yYyE�A�#��^��r����H���_N�ǌk�
S> �}.��j�E���:+2���eo�;��@�Z��iЧ�ɀ�E����hu�Z�"zHht~{kŊ��j�xh�A��5�ǇҜ>x �B�>�v�b���+�� {��U�|�Ð�vC��	b�v��9Z��se��CQc�I����/ґ���Y��+W��o���_�M|��*5e�7�n)Box߂�4yv*��g�,ߜ%���Êu$He��[!}+pkDK� %x[�8��n�2�9x�����~*���Ɛu'�/�C��h�������>%���)*�=��u��)օ������|���k���`cR���G�$Y�z���	ǔ��O�5ͳZ�{ٳ6�]-:(�gQ�Nm��mNHG(I
я�($3=����+J�)?�ܑ:�w��*���u��c�J����p2>�&3K�5�IdV�<��$�����nk]N��Wu��J�N�a����2�&�Y^+i�OY�z��V���a~�T�h��6��[b���f���n8����jZ�F�aW�|ro)�Ӻu��,9�� :h䈇�{C�#LC��W��B6�E�׎�nK�ng�����_�Љ�H��!2��س5{όL��h[��`;�¯-kkӝf3�D�[��'7A���KI&�YT��E%��P�L�
���8�(L�vz�3���{y�)�}T8�G"�#kd���0�gסKT[�˱������7�1R�B!Ɔ�ϓ�n� �# ��@V���m-��<�O���(O]�$�3�*.�>\E��ă�E$�̐�O��k�.4o.߇�ϴ�"���Tw�DUw%#w�b�أ�U	h�������&<��Jq쭃����}2
�jmjs;��"NG_&1�~�P4_��X���N����ٷ����5>��*���"
9�w{��
���9�ꖓ�i'���`K
�"n=�t7H�G��T�rL�T�Qj܅�TXn+�B���Z�콁$1n�3����T�D��!t�^�1�式k%;���ů�=@g􋞖��{�i6�%�&���A��9�r�+��y� xtUjE��TV|�e'Hy�߆a�7y�o�P����7���v����W,���K�Cȯ�)�)���&������t� �	�QvV�j������,Z�k��o¼�ny��&�:����n��PA�b����QeS�u�Z��^�^>���	i��f�K�+AA�֋�%ߘGN���yһUO�	a^���E�5�OT�
��~_ڑ�̡�/�E1������|��N��I	�?�DDX��ŏ�MG�q���/�O�� ʑΘ�}�P�L��Q�§4��R�r����j pG?���if�i��W��ݎ��Y�]㽖wʺ)n�虜�.���Z��#�.�d(V'@[0T��X�bMM =��8ݞq-���i�V���9�vڸķ��J�e�t��w�.�'I���MK���]�f�|����T�{�z	k���D��V�?U� [`#;^���⾽��u��&�V���ݛ��< X�h(���Ȝ�2P����Z�j]&b��#=�s1fyh�ʱ�Yd���/9��ǯ�v�b�Wڧ�F�JSǮJy}S�����{hL�Uh�R�ѕ-��/ �������?�J��P�'�)lQ�T�"D�$~$����gƇƈa�;���!��`���:�&� ��*��D��96I�&斧���I����������ο�K.EfZ$���/�*'�\ɀ1�?��������^���[���1�b�}ۍJU��*��Q�`m��IC$��Z[�*nK��I\>.Is��e����cw��5<�I����c�Yμ@� �<#���gVz.�|4�.�s �%"����[[����AޡƏ��{�Qۃ>^��#��j���ˬuryָgn��`*���' A��,$D�(O�`b��=%�L�V��rah'��"m8�R?{���>���]��˸�5�e5�)&GJ5�~��"�'��H#�H,�u���ǃ�{et�{�ͤ��dU�A�y�MwR��7��?�gl�M��gu~�8�\�[a�,3چK�v�y��*m�u��k�3����8�C�wl�B"h�麨���}/�yp�/���a�47_�4C``���O���m�ޡ�_��53�BdYQN+�L	hX�hQ6�D�{-��)���$_�Fh����7	A0�kx�ǎ,��3�L%��|3l�Y3}}�T��B���`��c�����y0}l�i�RM?M���x}Hy��u|r��c�H��!'��ù&���m#3"L�Bη
i��sZ��}z%�yR�g��(�J��u�
z�Z��eėu=:T��0���}�fQ�P�n�}�u��t�jc��ǰ�X�A�����z����oʥ5w�/	����u�|,����?J�EEA&Tb�NH��h�
)0㈽wF��M[��:�ܧ0dq�_�R���ߗcT&�b��˳}�Б ���c+ ��1�$
=$- ��{*
K<�6]|y�[�&B�h����}�3��{e���d��-$���P��7���L��0B�]z7�a:�qqβ�<;��5Ț07��Y4~�<Дם�l��Z���΀�@��";����x� K�C�}���f9��^(��Z拄_�3���%�x��oI
x��G�5�"�G����-(׵4yN;� o�a�������&q�å"�=�Э��=��u��F�QȞ?��~;�`?+M߬��bbU�$wLo�iˆ�Lu�\����� .tB��k�����T!��6&�H�ԳP�m�bg$ ݣ7����by6�k��>�o~�1_�]({���f�R��g���UO�؇���őT����6`Կ9�S�=�/�b�)�X�G;oU ����'AS�����B|�o��<>�(pRfG��m��j�c�fx�z/�������B���������I�Vk��wf�n�/ǃ<�	I6W��u"���ƙ��1��aZ��{a%���@�Y!&Di��k[�ڿx��<Z�*���B�j�tg%-�Cȧ�K)꬜��BI>tgޟ}�,7�=�hi{�	}x�7_��_�SLK^O�v��F��H"��� Ȍ	.F��AzV�\^Y����H%|O*,�� ��{�^\�O� �1M�mj-)�F9Ý��p�N�P���5�J�o"Z%L@�W����>?������0,�+���hQ��9��Y����[J�9C3��Zek�8��K1m��r�+{�~�����*]=�l!�!�zE%���A���Ӈ{��y�J�_A��M���Wp-8�����۳��PI��a#�&O�fwmW���+�io�tj%��MK*��x�&5����l�������}�j��{�@ӳ .�(w���l*�l��i23@� �¶՟�Rv�];5/Ե<ڗ%�NB�}�>뽪6٤���N�c{�\`J.v����B�6�0
IE�,ތ��V�E��)ڳJyN&��
H!�Z�X���6��>�}��G������rc�ꎠ"�kl�����<l5��`ƒS���0ƿ���u�^��j<�}/��M��Ob^�
h2�i<u�{7ne�|X=��3��e{�I�5g�K�4���kV`A8��h ��Ĉ�~��"�~WH ߰����C��i�k-�פ!Lh��6�;�wJEF8�������ߋe������A�\QW �O����0ϴ���}"Ca�
&��Z����x@�>	@m���d�S\NP7�K)%�0/zyx���N9�����{�s� ���k@.'.� (���3]O<C ��i(+Ϭߐ��L��+0�H
%�y�~���IF<Q�,� ys�)W\��<rⴈ�l�UEj\$#z)��H�I=u���d�!��Q�(�"���|��̞s(]��"�ʠ�6}��ަ�	��+c��u��:Ǌ*�5]�Ɗ���er���8 �d�i Wh�Au��=��9R=�?yL�D�״�iAݕ�*=���m�DC�z$Bͮ���]�&	��WYm���à�ٙx��D�B����꣊d��Xn{䊂����K�����^�6��h������ǥv�f?%@�[�#kl�-��)<]C|��3���}�="��k�D٨+�{�>�9�j�k�������р���S�ՏEI��Pcntd`�8�H���w>���Eb�S�N�M���ÐBI�zfq�19)���<0ɍ(��c(�I���"�����;�;��🪾��m�:� �����(�%$~����#����B ��K��|o���)��P���=�_��J�|zk�0���OH*��^�[�n��6�$���^�nDa�
;�X�t�Հ8�?d�a[RX��:�!8��B'��Ǎ�*Gv��n��Ҿ}�&��w/��,��n�.�4je��(�����/�����z����2obA��<bP)TM�+���老?M� �7.�e��pN"�ǢL��x�UP��0����,�'�w�O��F�7�䤢��췀7<
?��t=�v��F� ���d�̱R�?�u��Id��.�p)�����H���-��B�>�9���)0��!�G��Z��M�J. s�N.�bDq^��`)��E�?mhV^�Q-Zok>\I���;�Z�����rK���Q
l����_�!4��V#�$�S@�a�Ѷ�犊I��\p\gʹ�Oip]����j6T�+똡ЫMrb?�L��2\�������WY3�ɨ�+Ύ
{�����)���ٕg�%*�t?�ï�k��Gf��>"|��Pk�g�^O�s@3ĻWe�z�Uv��Iq<� ���'�1��V�z�^�$��
ڛ�G蕵�^��R�!d��A��p=��{G�=�������ln���6/�oT�����As�g�ͻ�~-�J_��}c��(0?�q��>Xie��cGD�!w���ۚ@���8=a�}�H:��pM��I )u�� TC6�#ٷ��qz���pC���}����1�Tg�g���)6{t+�3h�;��$�>ڣ3+��EzW�K�$0񍖤|�_M�5\[Y�d�!��%9{k<5��+�<������V6�x78��Rl�����er3 ׮���$�#�H&�Y�(F�pP�G]C�B/�ѫ����,E�TiIj�) p�>��.�m�i#��5�<�L���[��pNX��}�{u�j�2p��-��ƨ'��aC�����?�B����^
��:0F���\v����
��'v��ea�leEH�/Ϲ���ɪ�]�<������B�Ŵ�c�8��s@���:8�Z�W���vC0�y��DZ�N�"	�����G��g"O#��O:�X��à�x��v����l��2Q�� |u�|֣Eø����Q�^~�@Z�J�J@�G3�`˨,��ѵ���cO�|9�.J��Ah��i�f7�kθ#�x��֑o��,���,�~��c�����0�m�c��F�n�O�7̻�M��l�ʤ��@��iڹ;9§X��+��d�;6Qm����f�phD}omN���vM|Қ�:�&Xh�'��j#e����dڣ�<:� ��Ơ��
��N��oSC�
�iNg�2�I4hscI{��U[r��1�~�x�R�VB���47߱J��`<���|E_Q!��팒������6�r;vˢ�X	uU� ;"��ݺ�3��O����*��n�o�HZh��E"oF��w����K�@�ɚs�h�95��7}���p�Ԇt���78�ט�`'�+���m1Y����l,KIpX3U'�?��X[	��j�t��w�T�,'6&�FK�@т��M��x/�d�a�y�6h۲�"����a>W7���흺�
?"Z�0][�%���r����Q��6���`-��'l$�
�BE��>�c��>��	�e(�y_`�F(����C�����/�bUl8��r����t � ^���;ʺ�v3Q9i@)���I7E�p���T����$Q�о3e�T��� F	���XQ(4�k��LE�$O�P�@����v���R��m��xټ���)���Y��E�Q`�G��:8��!_ګ?�Q<��_n~q�Ųh���I�ؼ�I#��>
���yh^��n��-�$?�K!dMrӬ��;���F�G���ӄ~�)�*�����M�J����!���P19���_�ů$p�"i���#��mjt)�+M�n��#t���h�+��LƮ:� ��=�f>~q��Dx�3�a�J�����EGeÀ=ǽ�Q�s�S�VB�����xG�x�wKd�sA��{x�� cO�=I���<SC=3]�(���	�SNxF�lA@����Ҳ���,�29OH�lt�lQ�J-�5��8�H�΍AW,��_G��Q�n����T����	��[�')�M-�}�z��02��N�mW�[`WUEF2xU)+"�{���ߎg�%]��n�7ƢD�	%�\˲�>��i�߳�|5|��gOA��l$��$XM�r����H�C9�anx��jhaZ����`
��y>9��1Tx* !1b�(D_����;Jҙ�O���c �DL1�6T�b!>#!��=�s5�p?�tr��_b1�&'�y�n��ay���YS�1�ґWR�+��ӶoZ)e�4���}��g�G�~>�L�+���4�(�ɮӛ��/�L�
OI�8=�7/\
��e��uh0� ��f=ۻ�Z�}Ql޴�A2;�r�O���A��9��|�XO|A��ꀃ�S�G�8��1m�v;?у�[��d�0���[s��B�������uU��+g�u*gmptY��#)�l�#�s{s���KW�^�2�H�`�6�N�ki�r	�$������^�A�p����1�y�����#�xI5��B��Y%���}^?��U��G�K��)F�(��v[P �o5�@�{.@Q�����,�~%�����'}>W��6Z:W�?���Y@� E�@)���K`��H�����u���>Z}a��yl�����G޽k;<r�n�&uSI�)��hف,�.���
G&��U��
"�+�j�Z�����+D�V��Z�Ւ�?���G����fn�Uxo~�yw�Z��w�E��!X�ݶ��_�k�������Kd)��s����0~29��~��ƥ�d��1�?��H�����,+N/EV�;�2yoe+��薇���Qs�>�nI��E?VFY)�����R�}7���׬
r�޿t���i���݇�ꩶ���L��ќ�LX�>.R�W�¦�n��o�����*�ϗo�ЌZ�^@���'�#d���t�"��~��O�e�*����[�3��uv:��>��Z����],n.���\��_,���ye�f�6ng9 �:=<h�?�P��^(��vǿ��E��;XM��vWeYd(�ȶ�y�tE��Ჷ�Մ5���H�3��m���PO߅�/y���?�r�̝������6�W}��ґ�t]��
N+�E�Wm�>M���ѳ'9��{�WܱP���)�Z'�'��uA�y��
�`�����Pw�rc~���amԠ�����|�NA:�ĴL�X�`{��e�(k���N�R ���8�A����I��JP,k_R>�Ҷߴ@�V<��l?5�|�6�/Ӂ���.��2���j���!4��N7_�
�+<7'��ԇ�w惌���	2ڵ�cԋ��p7��(���҄��<t] �=������C�#��]������.��)|�6?���|�
��Xܥ�kDF%�q$a��6����`hϓ
���fHR�7Fq������$OP�Ő�e���k���?���;��h�ڰ�!�G#N�t�r�A��W�=X�a���ɑ��$�]а��ӹ^��/�(�� �(����K�����e.�|�_W0�Y=u��?>4ZQb�+���w�l���fqR9�������%[DK���ߊ����[N��4Xq�♖9���8���¡Qp�����ɮ�V�%��֟9��,їf[�[�9�͵Fs���!˙�E�$|7ԏ��c_�&�p�)�/V�z�S�}%�X�?�|%*O��Q������r:���"��U#���C�mi�&e#�.�$�J�z��o|>�D5]�W���e�������U:����~`��a�6���1;>;�	S#`��Gp�f��İ����U��SKP�p+��W��&�����_`�&n��`]��f�
m��i� bO���^w}����j�sè8�_��=5�
�9���	s�.64�OP��󰩷��)���������W�\
������á;��ac*/�Q"���L�`���-����y؂�g]C3���_I�؍Vx�{O�� e�A��,H����:S�M�g1+od��8m�^%���v��ny���d�vUKoW��&*�ܴsD���1dP�k˙[
��հ�������{$�����a��!�w��T+ �(������_ua;o����'N@Kb�Z�ؚ6Z��8K��X
��̙~���u�[3��%���TS�T{�/�M���Md/���b���B���RĻ�C�8� ����Hq�BaT�6:�����O*�T�����Q`%z;0B�W��q9H13�Z��@8M=��WE�!�����R�S/��֐��Bf�_����2��dF�)2}N�d��Qqg/
=��r��W��"0��ڼ���
KD�A��ҩJQ��b2E^�L��J֧�\qn�ܵC�U�~�F���s�pԙ��@DB���-���1�\/��e��Q��@&ۚѷ�k�Sw�#,���[�'6�r4X��>l\~2�4���֐z#EA�j[��`�G�р�$����ljgWNA&)�'�	�آHn��n�fK��9f���L��U���薲c���U�5_��n�
|9��ɨ�� >��k@''<�1��2�R�\��
@oZ�ފi��J�$q3Nj�q3b�
�*@@3��f���@Y(�B�j�����(J6D��-�Q�s̲#�z3�}I���6kѮםֺ��:"���n~`�q_�]mb\; ���7���,�.'<��Ȉ�����$��i��P��V�v��B}����ݒ�5��#������0@�gHL�Z�7����Tc]v�Ǧ\^������G���4Mx�m�syV�zY�ύ��&Ճ���b���N"28f'#6X!�6i��-W:�V�C[�ɑ���"�}��E��j�C��1���*�8}-�|d�4��Av#z!�7.����q�9p��l�ϱ�,��`*��KgC���*�j�&&�����U&8���;nM�vI�ߎ�=E	��S:�r"y�Y��ͱ04��a��ڣ>�u�N��3�����!M�pR��,��q��(S�?�V��U=7����N�Т�{|h�v\@����ynP�(���z���@�r��k����*�	�d���Z���F��C8�7�dNdge�W�20���`�;����xf�D�34#G�g�U;d�޴�"��������p�V�T��t����}�L0���!d{]���F�	���-�鶎����vE$\#��KO$��]t�Kbl�N����>]d,歠���b>		�G�7t�R��hiWu�����B~���G�{�U`��CkE�;��dXIz�`B��1�g}�T �<�W2�4&-�3=Ǻ���C���o�u�9f9�<�[Iy��S�=�\cւ�@02x�tSm�h����/R�J��ʺ��^ �x��;�EL"0�n��s��3���$��C�򬣸 :�9���h-�8W�S�Qb鵵{O�����:��x]��4`���ꓯ��P2����T]����@t�i:�~aw�f�ap "y¢9�j��8�����#
��p4��Aj6�;���D\7�PNN(����!��?��������
�ǭ�S<�D�����u�@1�ʎ?vg���JLn���h5�v���F���6�QXIZ�%�!2UhC>�,�
m�0Y0���76l?Λ����X��OG�|H���{�6+M��?x-7+r�a��H{���X�&M�^��"?����>Tɑ��\���}���L�������6G�B
��11�'Ȫ�$�1�~����cT�ݘ�1.���騡�`�(��joJ�à��R�?�l���ܾ;�3WO��W6�a��@Ht	t�۽BzW�7�.� �#z��m	�z��D{�����@;�3<�q^4-)��(#�S8�At|�P���޽��[���-m �d�r\�ε�TSr<q3��/ZJ˒o����a����yú__\v~�i��|��[�x[� �B4K�ɟ�@��¡5�>[�FI#���OI����ݒ,����&4Ɉ4���
qJ�>�@�y�Ё�SED$�>s3	R�P(�O�ŃJ�\-�����X)������[��\�Y2�/n�>�<[	=MŠV�K���s�������[����y#&{Z3�!�Tx.���C�*����#Sx�Ӧ��f~��U�[��Dհ�f�ʶ`bg���}P�B\��`y	x� ���tO��R�R?�#=�UN�WP@Ґ����V�D�m���~42�N/O0�xj��M?�+�����9���c묎3 ��ҝ�vP�eBKn�D�d�H��Z���n�wvx�=sY{f��|��m<S��8K������|��F.&��t�M?��;�X�/��;�����9�I�M�m�C)���q���X�2�	�)#����71�6�%x���a��œ�ksӯsJ����5��T��.���GEP7���A�X�	8ʬ�O��*]M)��7��kt[I���3�� Ml����9�q��li�i���i�J���<���*'[D�s���n�dE���Xȭnk_K�×��יo��?�7>���m$t
yZ� �^�J
X�4Â���s�p0�þU����ȳ�1��u��M�$��a�����a�8��V���pk��岭��cr�B�=�MZ�r��� a��氺�$��#+`%EY��TV��Rྺ�a�D��"c}��q�p�x�S��_�g�F9*�q۪W)=5�m~]8=��>�T��c�
�`Ϧ%���^ϊi�(s��|�ͱ�n� s"m���& ��i}WݵW��8T����#GZ�B%��A�;���һE� �+�J��KC���1i��s�>!�vlϮ����2�dN�����G�
Z����5F�O+uX>bh���Dhyp��r�������b���/�u�����B��" Y6 |�7C\�@dZ����`jW�P�X��6������R��_��aX��n�j�fI���W/��Q'��0TVp���z³\;�X�A��IZ��P)��?[��7r�I۰�KJ���l����f��ֺT��S�v��`W.Nx�����B��e��ݚ��>�2T儑s�#�挣����,S�R�26#�,����Lb�=����Л�i���7�����R���%�5��g6=L��s��$��b(��s#:b*`+���#��r�����7��uv<g�T	wQ`�p�ylV���*����FW�{�rGmu(��|��╲G!V{,��𩈡�ʎDL7�D��,g�
�ʍH,�X����m��çƼ������nTʈ��p��5
lݡ2�G�W]�/yv��a�_
V�����Er�di���GT��M�M�!/vs�p�L$	�JR����#gg%���LD��_���$�FuxH���x��aK�xA�~�qmd��Gk_k��Xv�����'.WAP���ΐ��\��B�o]��=�PL�����~P�|>>%��ep��"�Q�Xq"��F3�[;���dQ����.>>�Vj���&��1�G�<&+3g��,($��k"��uvo�F�{eH�
��A�5���̙A��X��U=k�U/O��R���}�7�ո��F踔u���8 i��H�K�b�S�y7��©�U]H��b}�M���n�ML%�q� 'Q��G੐���ֆ2����T�_R�ka&�,!��$C�������tC��D7E���Ы��A���qL�V6���A�S��(����
��Q""���+�Q֤T3� �r,��PnY�]K�ck7T��{6�+J��n�	"����������@8��#&e��O��[Q�,�`�Ha��R,Z�JͺQ�I�ߟ�vp؟gPw��7��^��Äm:��+��4��l1Қ=K�Â��g1���@t`�A)����7*֗�?�����l�L���ܬ�0�ʽ��z9�@��Y�|����x��X�����1gq���l��]��L��5S���>ip���\��*k-x�Ü��bza5�>�a?a�0�Ĉ�TY��Ϟ@��!ۧ�E5�=�M(��LHDD~,�M�M~e��������*^
u��QNP��"��&ש�\�m�g��OFGO>��Ҭ&���
M P��/����?޼��5�����AG�Hw�(����I�O}mޚ�$C��$P���w)_s�@��LnH���k��\�J'�Q���D́N㣤�a�$�/ͳ׃]鮃��Mo�Q���EX:nx���Ѡ�9��֎!:���#�!L&˽ (R��|OR	^�t���A9��aW��a�U_1�_ߜ_-V*~��w���=�-`L���1�;T�S�PxJՄ�SZ���$*,�7f���F<�<��r1Dx]d���c����7bܭ�;c�+2�!vIͥ��_�+��X!���I�Y<��[y�o-�8��H�����8k�q/��m����hY��/�rEY��z۝����^W9��܌Z�@�c�����e����M��L����~���ip�uGc=R� W�b���;�=�j�ۇVOY���!�}�4�}��?�eؾ�WH9�#->��"�q�ȱ�Ş�Y�^ղ%�)]�lc�U!-N%�I Q��F`c<M��D����1��B;R6��G5���(� �?,� ��,�R����Rx(6VL����
��%��it�>�Z����cW�#�#Fl�����b��p|��0���)�s���-��=<�vA���K���^Մ����֢��,��Hu�I2�k�k��E+��&����9=6w�[��>�c�$A��������.�Ey�a���#$P����3.�a@�(QfK�=PÌ�݀�x)�.N\5�v?�Ț�� ��Z���*='����IP_@h���H�/[��{�@��|��g��A����>,��7qc��=H�4W����
D#;r�q�-�g�����7�LD��w�<;Q�����Ϥ}�l����~J�c�XQ��0�X�с�!g�P)�ԅ*o�ƣ��v3��E5�v�����?�#P�_A @RƁ�.��ZF����B_'���X�p�E#ER�XvUNb�R�2i�ݮQ\�_�Zl����)�g!�	H��o�ѵ��D�Vc����w��Ǘ)5�h4�D,��C
�$sR���ފ��5�%�mU%f���d`b�Rt�71�gۗr�﷐��!t� �q�+,d�-��=�+}��4���
�>o�c�)��?DIg!7>^\DD/��`�`m�ܕg�>r��E���^���c�ua�,v;'�rY��K(��
�4�掵�7�Ѵ��@f�&��9㦍l��ӓ,��j�!�#�hh�:�܀�œn�$��������fH�d�>��3 Z�?�i��Y�j4E���08���_cI����k�8g�a�����8���vZ(H�:�i��{�bH:o�r�a+�7���ב���]����-��_y����@ge�A���)��$\RJr��P�9(����o�$=���\��^�q�֗?AA>���IB:�n����(��ָ~{�}B� ��0�����m�ٳ�d#@��G� g��d������ʝ��h��-�����$���Q\��$����lW���m|h᥵�=�a���$)�H>)�����#K7�V��#��� L�k�H;�r��Ǩ.�3��,d��Z����&�#��,��/S�%�Gy�X,�����p��𺯯n�:3~����`��Ɏ#��I'굪���l�j�(��&�J���t�X��B�*Ot���o!�<�JH�%���hW;��;���Vۏz��M�ꝼD#'�?������ ��u5�0QC�3X��_��'�[Ø��	�N4O!�3�Q9Ҏ ���G�~h4��M����x�p��h��b�-����4�j ����}�+ĳ�#��7s*�tX�T�)׳�I�œ{N��෷���y�q�^K��po��S�ʗuq���7T@����$�3�.���1�*���"��f�WAh7��8���k���wŬ�V2g����s�q;���z���!6Sî��&���!�[F���2i���������6�9�ڬ�~د��led�t��D��P��kO}�N(W�c� ����#�_���>�g#l A,c�M�A4����i��xeA~�tÿ���
�1{��!l�,�y�_�����[�>
�F��Ν�LP�9��3W��������;���ۛjeޖQ����9֗��]��X�oj����JI���.k\�9��:�޺T��M�NI��s��+W�J��9��+��ˑ��% N:V���>����T�x}j��#qE.-����e+k5t���tߡ�GgO��-���W-������C�����+�`����v���9y�cEY����f}���YLR��� ���KI�����5.�y�њ��[V���ؓ`�nw�|yT;�yy"Xa���%2T�m%�	լ�ضq���G�B��p0�������00���H��P�X	:+�&��-V'#�L�}L���{?C�C��}��>mC\���l\�O�F�ƶb��A �Se-�ۖ�a���3,b���:��k�`�Y�a�gF }�S�܂p��W�Z��8�,�Ol8�@��	�練�����T��|9Z��RП-
�/��C����7)km��+JH4Nd.6�	 G}���6a}�Ѓ5|c:sL�'6fٿ�>�R��1�D����x� G�D,E
���tZio�=���9��IV� C�ph5c�o;�b�B��'�� 刯N��'���:�� ��+#�R���N�H��1)��y��?{����p� ��hyX�(�6��	j���ڞ�Z�'��c/n"�ߞ8�L�hDx9�Z n[ތ�(�t�4���ǽҡ%Χ�����Y͢u7��}�\t�N^բ��e<����j���rk	��1h��3�����i�CM���ǿ>�q��QE��/][Va�'"��i����tf�c��O?��
)���U0���\��Y��kP�Z5G�6����è?�ck+�d�{QȻ���hI.{�q"X�dꚈ(�*�_KE���;�!�Ŝ9�/�d#�2{V���oΦ	�c����,��+&��z�cN= *e\���K�MY0��¯�zդ���q+y�jo;�#=�R�D�M�J�(��߾g�,萼=c��ʮjSɁՉ��U�|[����?�&`_��w��ɵ�H���>%fgf��	�U��#��[�b�9�Z�@�z�Ÿ%�`#p�r� �+���(�P0k��]��#	xg.?����<��R��i0����+�h���kD�L.�<3��
a@�?"]co6z��Q("����}#pz�g��F"����:��&1g=�"��M{�A -1*;T	J}:��
��ΞmѺ4!�*ݴy��;�4���)+� ;��aFiw��2�����69�$>����Ȟs�6� ��b�G���{�Y��9<fW��_�.����kŷL�E��t��Lآa;�`�[W��Y�d�ѳ؊ܵTz����@���9*��ު�f1M��s�w�����D=�Lw:���q�F��A��ScH!�FP����O9���g�����~(؛j�L
��2jK������#�8�J=X�R�x7�-�S4��Y|��nI\"綨?U���5X)ѼoXH��9k�:g�}u�A��M)��梎��mC=W���-�~6M�O��
�	]���lv&dMs�y/s����ᵶ�ة���D"ߺv�j�1r�p-%�3�(g�{���8G_���5��J%:��Ѽ�vz�=��t��2ᇎ�/ B(-bb� ���=PY��yƘ��⅖��eca�B�2�d�����i���|-n���ߊ9�*j/�c�Ww&��*�4�G���]��6�b�;F��3c�s�Z�DI��D<{��~��5ݯ��Q�7�,U�9v^1|B�ow�����|z�,&�b��7i|�U�Ш���ZA*���T�٪�_k�.[���8%�)gk�ʬ����#�)4��)�V����ݨ�a��:^J?��#�h��時i��\��Ȼ_P�� uv�3(�ݚ
���֮5�,�GX#�zQ�Y����I��#���FĐ��W�s�&i6��%���Ͷȯ������ш�B.�m8������2��>j>LSʅl�s��Y~e�0z�}��L��&�6�c��٩�aW�ѧ~����G�E����v��脰Ѓ�����>��B�fٳl�MfW��lm#"��~�����HD�WR.��s��ܓ4v#�};��ƀ�)�q�������Rb�q�5a<����p�m���v9���Sh�Ȳ��+ �J�+�=o"Յ�G��"B���"���Y'�iܗ�%u�/nf	#߂��Z���Z�#e��R�;Ad(��L	1����6����y���ꦰ%�'���Ģ�7/\��������P�/�L2�Ѷ�8��t�#���+!��0�S��sTf*星�7?�[��e����	���>k�&���c��ʉ���]�+���J�(;��b�����@#�i�yPIo�՛f����{����<;�ү�����"���עȄ���x��k=gJ�z5��4�=��(����1f�ƻ�2C�I��[7��S<T��X�]��2~;�0��ˢP��XJI�3^�ř�K$lJ� Ĩ�T�@�lO�I}p1�:�8�2ۉ;,��Cs]%�}Qf��Pߋ�}���>�dM8{�a��_�h�
���L>9�M��`�MSШ#�*j�d�Y�f��(�]z�Y�PC7�sߗn�)���K����R��
���:��bA��Lua� W�.�Qj�S�pQ<����:d-��-!�w�F���]���� �]�!�#A�6B�2�ޟ��,��?��h,�B�}ݯ׾'�N�����@�lZ��C�$a�pN�=�����{��;0nlc6�/�/��h��s�$Q���^.B�NLt
���y�4L��|Wfgb���kۍ�w�%�DW6�R]=Ѐ]�8��8SF��"�$��I�0_°�q���$��H�XJ�]`k���nV�p�D��y͛%�M�������~�;>I���5̾�Z�OP�����"Пz;����٬����E��S5[�|�>�k��r5I���k.�R���<�0��s��#h�ڽ<|�L���f��^��Q�
�K����Ѳ��c=GT/��f���b�&E<�ׯ�����ay�Q�[P���6l����h^T���k� 3�|�r���߱93Qєw���FՔo��	S�j���HW�G����K���	��6~5�������H)Gh�Ad���;A,z��zL451��v�������l���N�ZE,�A0��%NK���s,0��ޞ�ɕ˞����ًa=�� �l�+��g�tp���[���x@T��������Tu|�I�Լ:�o;V���n�a�����F6)����IG~sN���C�<��q5 �sݧ��]}�gAt��?�J�h�<TA4\����9!��L1�'m�@�S�+,e1�N6D5.��SW��`Fv7YR��A>�}��]a��	��*�}�1W�)��	JA�_�L�6)�>���W7���.J7�a��`I���w���]�NM�5/���Z=�������<����EO�����S�A�搨ۻ�ו��9b�Q��@/r���2�Y����|��G���=(��҉2�H��F�C�$�|�Os�H����S���i�ҡ*z�BsM�S�O��aʍ���ޘ4-%+�F.�+x�r��[$b���p�����$atZV	�H9-�����D�@�ym�75X�<���ӣ��[*c�?�)�1�	p�����_}d�jW�߶b"�U���8k��'�p&�M���Μ����1�/
2������'�����=?K�.g�Y:[&�iZ�Z����s��ݣ��b��q�Fb$�(Q��e� ̽!��ep]���5���t��#mt����`��V�P��	X�,P}���f���l�1�)#� �l����U0�ع%,�R,�V�'�П�>@��c�W[�a�,y�8�Y䗹(���͂]�.��F�����.�o�0���Y*�߁�$��n����� ��e{�]�O��|
�~��Ǧ�wW7�H�43�9!��c��=ܒe����m�m�>���ޑ?ͿBD~+ͥ��8q`q\��j��m��xx(�"��?֊1�S*p7g�'�a Zr�z��]��C�1 `&l2�'H� /ku�t�w�fK$�+��O�?9W��B�,x�z��&u������ ��k���}׺�HZ�MY�'�ڒ9�������(� Se�c�Q���Q�sŋ�-�0;7b�Y��ܕml=�Q�]�l�-��`.	bl"�7��,�v�Uz�	�ݟx���ZI�&�MՋ֥���"R�^ď�>Һ��	Sf��������6�M���#�V�1�T��\�Fo{���:�R�;Ȍ{:������ڊPt "0����3�QM��oޱ���c�z�~���z��jf����5���y>Z��¦��DA��}�<އ%�
	���;L[��H<#�'�;�qu	��� ��}���#R��t&���}5�E��i��"�#�>İ���	����ODO�m���:���Hr���.���]�(�$�f�:��C��A��e��0����«U�Po�y0 q�ʖ��˘���)O���m�v���l�D�O$мZ5��9p�	mW�t�;B)��(H�c����S�#�kj=��N�ч@I���:w\8|9��hì�tIRx�L��~:��#>��(02��]|[�ǥ��k��Y/�2R����}���a���b04L�FJ7w�)�ӓ�1b�(��2Uq�Nu�f��/�-��9��C'�o�=x��$��w81�ƑG�s�����5P�2 '�怵����s�e8dXY�9��c,��/���ņ�����PX�^��wwm�hO�/��K$_ʠ���`<����[�vHgJx�q
|���Ii����2�}%"��bR@U����{~�\�PxJ� �#� 0\�]�=��S:���c�p�m��otXYz�D��q�?�0/)}.��_zl�B������>����+��薋�C���62�.ܻU��t���� ���,4~<��'͊��H,�&�2�Rj�;,3��vYb�T7�~8$w��,��
��ػ�)(�gNz��%���f{d�xki�]���缍=�Mb�~U���S\}��yޗp����!��y���/�r)���|�$�	���2n��_��w�����/���/�N/V�>����w�~��rU}$��	נ�4 X�{�Ov-����玕ß�8��ʚ��Q�*�U�u����	R����o!��Pn�F�Q9H��Y/������4�n���I�B�&�M���i����z�����ɡ0�7l"*	����Ћ#eg�1��r��?cߺP���/
G�~��<di�'�	ꑁ����ل�y4˘	�%H�8��O�)�*���g��|;���:l�t��z��nh��xxg�|�M)�AҖ`�p ��A7$˜���b?8�.����&=�~�y�Q{ో�%{��� r1����Z��� ��##�J7Mز�zSm�u�~t�w�����^�aZ6���C�e[������-� 4k��K��V��{�+B����CҰ�cfx�q׮�Ul�ţ*��o/\�ފ�t���"!;pa�P͓�}G&�`i�2JPTSW�4�U��^w�Xwn�?7��^ߌ $�%�|�,N�����uO�t"/g��̠����ZS6�'���k����Y�[�����w1�+�3�����N���0�&|��'�	/��+bu%��a�B#r�ӧ�l��,���WS�o��N����j?��r�`���an���8CEt��z�����y*͒�z��Őc���<�57��p���y�4:z q4����Z����]���`��$r�>�G=�;~�{�������G�
4V��T�x�C�	ݨ��D}��N��%���t�R*����T��/���](/rD�E��KB��=:|A?*^��3���$����C.}��kץqF ؿB�BDj����m�_h�
I����%OB��p5	8��T�&.�#��9̘��Ӄ��V���ʕ��ک������V��F4!!��_c���!�T��}�<j�a߯�\w���c{J�M�x�c�"�F'�JN"
6��2�X<jc�Z(Lՙ�iG��։G.7�  9�cS<
-�[���D�E�*7C2���@�`�Mc�Fl�=%Z_q��;d�柰��"������<�!��G���N��, Q�>t���=ì��&�)F�r�U���~���s��|�h�8D�ϫ��s�F����\��>Xd��~R�s��<?�i|?�n�����?�j`�ĥ��a��K�G3���N*ZF�qb���1�mf ^��ٖ�?��j�L�H�n���^��
(%0��Ɒ�����!⸢�x��'�2�����u�kL8����xҵs��K�H+J��Z^^`8���j����������.�F��Lt3��1�ݺ�V���n�wr
�Ϯ\%S�p[���o>�Wv?k�θ1gE����?C��P4�
I��6�����ڭ�g[�k�'��l=oRc,Y;�S-��5x���7�p���g���(�B=2�%��-�׈�ees�Op�,���̋�k`����&�aZ+��R����}:�����h�5��T�y%�Sfb�[�*{�G����j(�9r�M�H�'��U�@	|�'�9)9��;�{䁥� �Gv��T���k@ę�4I� ����q�K�����҄+�T������'�<8K�a�����6΄��xs30�J�x��Ѿ�i&�Ŭ�����k����a
�a����o�$	q�*3V�r�~e�����aNK ��%&~Ib}5N ��{�S�l!�rY���F��-�D�,�����)�1��nⱟy����3��
����Ii���3�qlu�����΍�>E��m���g�b
F{b}����8��{5�6W��c�o����/g�g�~x��A�|�*p�<�����zq��4��L*���gE&g����x�gAJ|�#�,e��Q*>�'�ݥ���BM5ܟ�W�z�r��	%;�i�tZ*5�����W��ί%b �j)�gE%��D� Stz/^>3�9	5�����M��>lBvd�Q��[�,ݤ�a�Eݙ��-�9*����G����n(GyeMV�\�"�Q/[�3̬>pC���r�@�>D�J+���3E$�g��r�(}K�-t+�Q4y��F�*vţ�G�o�vA��┉9u���E��wB����ѿ�+;��A�>�a�Fz�Ғ�x���D`	_S�������5�K,�[C�X�M��J�y���-&|�r�u�>h�V݃�������Q�,����+Բ����Q.qB����٬Od��M�8�y���ߍ�Xa̫�ֻ��-�]*�訮���AR�Y��I�,�n�b���4Ops��i5Ef�F���R�ӭn�\/�Ƨs�g(I��zd��0�J����/n�=��a��ty
��q��Fs�d���S���[툥�˝@Q"��{$���h��`�aTD��S�?X��M��]i��.�Rڇ�G�ڇ66���ű�e1���f��vZ����i��  �`�����a���X��:�Edq\gHe��.ɰ����1����l��ꂖ �`�&+�1Lf����0�
��nkv3Q��s�|ù�5]8�e6"���pBꦘ�qD��CE$�7��{\�p�U�I_��XL�y,��'E�4<��=��D�k�~��}���/=x����s��]�tl�g�f�;�n3�<�qm��$ct3��P�����A�2 S�e��V�s[@�S�C"s��:Μ���;/�8��A��sq�(�v����&��4E�$#��Ψl���|��	ݭ��7
��f����aҪ*���յS��S��=�r���������C��ӂghtѢ��q�yJ��M�?���<B����&.��A�S����F^�з]�^�E
���\;��zŰ���蘵���h����Z�ķ=(5u�g},���hb�i�����g!��Vi������Fp����:��<�*h>�UI��Pv����x�͊1��5����e�zw��6�Kqe�Y�
�oڦ�8}�c~ɂx3�Qŝ�̹(����l
t��=LEG�l3Zԩ�-c�Y%j��X�u~��ٻ;��h�����l� ��Ex�T��0��0���1��j��:_�<@z�NRfꋮk5��;Iľ���p�����n���&^U����;�J,�.s��rX�qG~�C����$'ǭ�u >���Y�p�fJ��Q�{���`KR�_;?�?шf�Z ���?mL5,���Y1G���uTAl0�������yW�'1�Ć|��r+���k|�r��XM��v���#����y<y�Q	X�
�R5�A��T(���nض��#*[1���/��Ӕ� *e&q��W���~+0ny��+����3f��"�3M�Ȗ�o@��\�|c<�k�mcD�χDa��p>]T��A,��u��
�q�Z��Lz5�&�/�&`H<[��)�2�k�9�K�?�H�*�i�jj�l��[�����yZ���Xn����-�]���V��rF�5.o�ֽ[�n	����ԙS#A���d��؏ͯ%|��_*{�\�b��}gh3����ʸP�O`5u����י����4L!�e�6�A��p���˥ v���{���2�H�����@�Q]�Y�A�3d��?��ᣬ�����|��T�*�r�U�	�؝4�K�촙��{`��`���U����
���(G��߰�`쏂�OyO��_!�v�#h�<��=ԫ���Ȟ�$��2�p �S��B9�\��%�"+r/m7J:oޥ-z��@Oʒ
\����V�o뵍3�cp�S�d�)t��8�d%���ml�o2|qT멠TMŰ?D{�n����gkx�rg
��
HHz����a����z<7��`�=�Dg�ТY���1��W�oKZ$��y~fQ_1���{�:U~�O{�����5M֫��'���a4�w�O�
�8z&��Du2=B�]%� �jJ��WR�n�:ᣔ�!�:��-����Ş�LN��U붰6�����6^��%4�֕�"!�Gy���wD�p6c@�3�y\���s%˖L)q�����l�b3i#��<�ʺ,��Y/G�i�Ut�����P%^_�S&b����Γ��{�TX�R۬bsX�Hؑ!`��gx�� ��^	v�J"`VT!~�C����L�ۆ�����}rw���]k+�2��i�(��2��-P��K�ƄY�K[�,Z0u�]Bf��:XWm�`�a	�ݺ飣�x,ӄ�N�I$U@b�9����W�%p��j�z`���H|
�B��H�u(�.m=�8^Ԗ��O=�С�.��h��9�w*���߸�f�Nx�8�7=������5+AJ��B�����׵vp��s�*ᙛ��!��õ[��[����4�}>;ɲ��QA���_21L�������������
�Zi��-$�X�_��k�ѱ���U�ධBwX�V�ci, ���w&������/�Ҕ	��Ҟ���ԛ\�����Ê.���`IxVFW�M����0�b	B�W��8nF����8hnj1Ȱ�S�h*W3G�������)4��J1�m����@�lL_��n�l,z����|���Qe��e:��G�������γ2?��K�n]4� �Y��Q�*�!�`NZ�Y�����*j��=�%M�6s`���Ҕ*�1//�}��+�Ed�V��d)���r��Qv�H�K^�	Dlh�d��S�D�]�{W^_@�Gw�㵨��Ŷ�"�س��h04Ш2M���f;��ݤ��7��q��p%��D�H|E�^�E����Օ�c�;�����j��B9˅#(���eH$4��C��������6ԏ�}ں��d���	X�l��.����G$��Z��͑;����=Y��K_�lBZhs��Y���@P~�p�A����cn��(6w;�������>_���[�\���"�Ƥ�+bS9!ӯ�F�"Ō��������۷��=oӃ��@�1�Z̐ٓ�:��ѮY�O*I'X=�)�i�;/o�[���UػV�&�7�ש)-�綍hQ��D|����	ӥ2A�12����8��8���ُ�_�{)j�,w4��k	��D��e��jl�<lZp���Ȅsظ7?�]�q�dx�ֵ5���`)rsS����[`&d�L\|�)�b��;+ ��ۤ�:ʶ��� ������)��L�Ȫ���52�y��ng�
j^��1ۣ>���.����u��Y�($vW$|N|���6O�?�(ɦ�����Ei(��y�*���B�����; 9r�����@W���>G1��zZ�͞��Z��	^:X3.Rc+���]x��S�P ��O~�2C�!��*��R?;��% ��j�}FCw���)����9�J+}Ue�H1��$���B[��z�L������@�3���^��l�m	��°��<�5����[aM�
�^����0bMދ�ګ-M�^���&��ҺTȷ���[N�E�D۹ղ��b��]V�
�:ڦ��U�`���|zd�h�C��_���;�'���� ��
�}��x]}=Jjх}m�,�X`�٣�Tb�}8�3	�&["h}���u���Q'zAa�tJ�����{8�[�Z�y���%�gx��c1����Y�F�Sٖت�$/���W��;�Ug�0N�����G���q��� �(�IF����5��P������;{���������Y,:�*�L]d5�_�qq�y�<Cv9�$ypľg���� �ӄx��z<T� \
s-ˠ�z��z|�:�.��+��b�Q(N�,�ؠ:��!{|�[��]�S�q�xO�MvG��M�DW.�i��<����R��a2��l\��@���e��zt� A�Ms3�ՐRm��@�yJ�i�SXZ�/���7≼�X��ÏPP���gqZا_�c>��	�K@�`Ҁ/n*��M�|cǤ�W�^�4�깕|X܎`�?�/X4���,� k�$���۽���ɝ�V2��6rX�xw�`�3�k��e`k�M����`�h�k��-��	����Z�,����O�u/*�����0M���Y�}#��5{i�� 3'&r�>`Ž�u�g[k ~%��fN��.�4H.2�[�1,U�O�L�ka�t�e$ܹW��P�*��o]d�;¡)��j�p����b�mGMۙf`HH<��W�oG�D�1��1�O[�̉�y�
.�G�U�ӁEZ%vS�Aw�98�?���l�aE6m�g���:yqyk~jr�hް,��eڷ#���ױ��W������+�ߥ�u�ur�c�L�~L�f:`�A����"���/m���y��ɠ�6Y�˹��S���u߭���s��i�;����� �Zb}}�"fZ;ρs�����x�60�n��~ ���& �"��4ӱv�;����T��e�������$D���2��H��![���0Wn��ꌅ�+�ۅ��O���ct �p�����Oھ!&(�-wrC�z����q�Ud|��*-U���EI�.��5d���$7:�È$:A�M`���� `_чN��|�u�����3�u�������H���w	]�n��WS��KC�,S���PA���)MQ)������!ʍ���1'�#�GL��6l9(�)��㋸��p9�O��"�"���������_Gf嶃.*P��U<��Pq��گn�r#� c�M�~�l���1�B�,*5�����<>Lvj��^c-h��$�0	����3~�ퟡ'���"����[��-OLb�A�֤�3YM���0�M{������LU42D6[�`����}G�N�CT'��#����[	�7����α4�җ!��Z�4#���-qSaCqt�������'铃�Զ������ғc���W�l��p"����?�QL- ~�8W���F@��a�)Ό2z�1�kr�n�+� wG��*?kgh4e���T��T�e��S�-s�[A��ʚ�?�3�����#�L�Q�V���G���1�،&':o����A�����4������ʵ�b�~��u�C�o�=2@y�������t��|W�O�����M(���v��2�C`2kxP����(�����Q4��4-��H"tjs��K����+Z�pA���V��u�: t��B1��\.����5]��h����9կ�24�P
Fh#-�G�gCQ���s�|1�E��O@��@�h8W�"{�����ڠw����R�������:eS��A+�)ѫu�]y�{:(���4oQj�0��Y���:��S�O������y�b҄��D�b����C$稰~�B��j�m�)g�X�+�!�<�0K�E�x��-Ot��="�y�JZ��xw m��`�\ϭʜ���e:��Eu1M���)"X��M��7��.�+*r����z^�d��B{��3)�go�����ᶹN�r}d_ø��(w̓�3p�����V���آדnu/��p��|�$��29nv��=U���Mm�Ǜ��s��4�q����HW���7�}]�:����j��P/u,X���΃؉���nm�3�w�����e��XR��J��;ES�������&�01��Y8��O����7E���A��S]���ֱ�?�n����7�W��w����^̨My�&�k+��.a�#m��������K
�침x��l3]7wxE,�b���0����/�{�.��M����������(ٷ�!!B��]k�@��0��V{z@=�$DA�>��U����?�nF����Z�(6ߠ��/�r#���������Q� �!un��ۯ�_^���ŏ@|Z��SeT��k�F6i�[�E|]��!�z�-��M��LǾ+l0\l	\����6�&�M����,glţ�t�X?>�zG�I�]��SC��c�X�Y\k4�6D9X�ڋ�n�_l�v��D�1�0OYe����ֵ#��|��秬�	6]nO��0_H֛؅��Y˚:"xi�p, �tuQ���� �� ؓ����=0k�{�4ӽK ^�ʫ�l�Lt D=�$}y��vp�R�R�*묨�%D���G l"����~�/ϔ�2Q��8�B~T}�Wv}���6����0)�Ĩ�,��)��y��( q��x�arR�ϒ�~�rN2�Zq�U��K���ǻ�tj���2��ې�!e��i(d��@v}#�T�"G�kPx��*&���(�o�88�`�o=Z�+��9׳#K*&��� T!/;��I:����!�&|Yu��G���>R��:D�:�W��Z�"vϽ��ѵ8�~�6k������h:�FF�惬�)��on�q�m�IZl��J�C�
��Nhׇ����j��U�ɭy�n��ҵ��۔���~D
)5����Ǎ��tng�JRU�����\��9�7�%�B5Nһ9V_�
�j\3�Z��;P�����Ș�mY֠͠���M�I'F����XtI	=�Х�j-6��!Νӫ\�9��u�0��.���5H0��zǻ�I_'��5P�FA]��JN�ʹd�����P]~��sR��7�fb������z�&t���R��>O�{���3��E���po0��7������pcir�q��M��(�	�\�fҼ����P�ɲ��j��٤#�g�`
B0�35�ǳ����QH2uݽ�n�S �3�]%L�N>	��Є֢ϥk����פn6V¡�7��"i���[�F��=�b�/]f��K���5o/�o/H,_��=ӑ_<}B������('>��p�8�i��8�GZ����E �m���V�����һ����a�G����+�6�BO�=��Y.�K�Ʋ�J|��ud�J�٣M���U~�,���m��fѮ�30f2
Bg�3��0�K[�Ɋ��O�]=��VfFl~R���ܻ3�y�ע����n̦�#:��yE�<o��n��ѲQ�og�O�_����*�p�b�����Z�v������8^�@\@q+'CX$�G\�sIǸ��o�3X���ER�X�(r���WH!q�l�)�:ٿ����:9��s�S�W��K�!*^��M�`e:�q|^�j�j�G�}a�lh��D�<�׌ۆ��+Mjٯe8�WK�k�sN3� ��V=�|���VD����\�A���zP�����-'��
�r�ȟ�Ɲ�;�]N�7�nE�
�c;!a��e��|�b�_�&oi�gO�G�cʏ��o������˿��j�][�0�d�Ҏ�#���
�p�Kȹ�V�^`S�Z��:��&d2��uII��yy���|��V�Pk����'��pq(�>xC�r��I���ܴ�����p	�9o���\q��m�]����*:���~Y���d��I��6�V��-{:�"�L»𤩓��^�X����ߕVUaFpB�O`i��M�.0!Y��s(���>�`����~�q_��v�@�GEz#
	á�ZT�@(0P�\�9 ��� H�����м��A�/��:����_�7���	P�5��P�|$H�1or.
���'0���p��D���HwUW���;��H�if6Jf��蒉2���#����"B�#H�f'��\����P-'.�آ �I ��~xȚv�^a`G��jk����;���~�v���.�J0�O�����H�@��)WG\*���q*<��r�Z�7�(�=��8v�i����B�c��&�
��&9�~�
n�[wTQ~�_B����M�P�L��Q'�U+���b���;���ɲ��ݸΝ��y��JQ����f���W"Qn�3���Ľ�q�q=M6�L� [nI��G��
ѣ�ٵ7���#Npw������:�Yp�Jp��r]~��z���p.���� P�}�"�Y�|֬��y� zz|vS�e�^dԽ�`ҝ�
e07c��]���p�����֋@\w������Q�w�o��狍�xF�JYP� ���}S%̭���d��E^����}��:�8���E)���؛<��7�2L��!��2�wy��!�˂R�s�8ݩ��Hz�m��f��޼���*F=��0�<���5���ľ�=o���?�T��E�*]鱲b@\��E1`�YU@I� �c�+����+��gn_J���!J�R�o�;@�Y9��+{yc��_T�/��L��~����g�*�����A�w٦V���m�Q� �Ȁmv��4^ԩr�VG�)�x�I!����U�����V��2�����V���p����4��� /2	,+�Z�7y~}Cj�8��\�rvO��VN;��}���;Nu/�;#b���R��M���
܍	�1G!��j@��FK��Jea��gm՘O�k:��U�i�G�2�wQZ2���7?&X��9İ5�`\$U#�pӧh���X���";�F���J;�]�iX�|x�j��,�`�7Ȟaof�T��\��փ���ի��8�	���y�����"
`!���S�Df��s.rU�q��l��6�W1�l˲��)1��$W-3�DU��wH�؟r�B��Y@��l-��y�Y�}Cƨ�N��=��#t��P'O���E�����KR�-�J\Q�Zv8�BE:��%<9j*4��$Q�ήvwg2s!�UA92�P���o�b����VT�����tV|�g�|5����썢���"�+�t�זQ��rZ�3l
�J��b�Ԭ�sH�f�Q�}xj��ɹ�����!�ǎC�S�q3#��N\������o�OV�c��zwO�#~��v�7`�Ի��@��lN�4[`֊+`����P�b֟$����Py[�4�Fttnm\;;�PAX�j1�5gmq�/
�~ƈ ��J��P4r�D��˷����힥e��]M#=���%�	�?������8���ylde��T�:���*����k���Sm�?��Gv�"�M���& Ĩ�����3} �C�7N�Rl~c���5�<�zf$u�H-�n�6}���	Q�^�W��zr���ɞ�zx��B[����(� �'��ߖ<�l�L�R������4Uq�}V�&{�,%-���S/���l��[�)zȘ�y`ne�TR��D�'�0\;���W�F������߆��x\ (K���V�AޛewOS�W��>^B1:��5�b|��iON�#IoƗ�p�5[!�����>[��C�* pc_|�28	��Q!sM�A�u7U%"��p?v3֩�$�'��LY�E�8�O���c;tm4���I��s�#�}$����Q��
O���ݹZ �o}��^�����{��KK��_��~R��(k�'af������O(�蜂q@���� 4�}K����8O2ņԝtM?�W�����F��=E�F���>e�|]�O��Po�a�v$��cSj-5��� �r��9{�x���Q`h����,�a�4�F�l�ʍ��.��x�%Ϫ��ˁ'IQ&�{K�T�0)ځd��!������ ������x/g�!\�p5�����S_��.:�j�K�+��I�9yN��a���&�s��s�V�ˌ�S.�jHi�#~���;6�wͮ�U�q��-G��z�ho1�)J����6��Q-�r�F���*HY�(Q/�M�Z;>���6�$|�����l��5�bx2�5�61�wi"r��V�ؑ��j�1�)��ܣ7Pt�����k�x�D�?�0g~<rw�DV�b^Zt�}���~b^�$_J�ay��f�=S�Pz��3�*3T�&��~�u�Ϛ�NA�����-0��sa�Bؿ����ć�_hݛ�Б�F�C`�n��Qś�̩u��P�����[�Ԝ&M��_��֢�mgf#���M�rC�D ey(⓻�g���RɁH�����#�ҼҪ�]H/,���@�<U��+��1PDGǳ�U�Nx4�Co��l#M��l\m�����V�hf��q90�e4|����,���f�z��aLx��B�Ƣκ=t�P�6e`)�;�� K�O(��T��ci�ʑ��nl�eR���r	��'n���"Lz�V���<H�+Q��{�ʬٶ?�g�ߚr��+�������[/.��66��-x�	z��8}��q���&��H�ꀕ�~�+|S��k�|�>�<f�+`p��%�6��A��5Z��k��D�������1Sk���r�9��[iܩnA>�Ū3�M��`�|f��1�hk&���m������Ob���0�k X�b���D��.@fw����[��` ��6whV�t�4F
֬}o�|��4�i�ã���J'ZA}m:p"��v��T���U�������j�]���F������}�7_�=�rE@L*�{�32�r�$� o���w� �gܬ{�.�<� �E�e�G�]j!�eB|�:��/��tE����h�-����E3H�Vv/�P�L����i���������,��d�E��H.ܺkh�3�jW\F���c�m5���q<�v��ɦ��ġ�����jU%u�x�_c�X�,G~B�6'��-�#| ډk70|X�ɫ����':/��c��`)6sN,���]�Vו��]p�Pch&��E�^�X����Y͘��(y�wr>�g����\3*0�Ȯ&[�cVC�9�F���� i7��@x
�:{�??�3��t�8n_6�;5Egf��c[��٘�α��V@B�i]}����Y!�R2�M�H�M	�*W籓qĚ����/�r�:�q�<cn ��O�A�D��_�Z�ʓw ���>H|}t&���mz_�!#���O��98����(���ȣX��8��<��--u���K(��~��dQ��E�� y��434����˲�ҵJ��~g�w�\�����\{�O��
X���#������c��~���>�$����>y���߇�e	r���g���ֲm���V����ߠ���{�Ę٫ˌR�4�CS���?��0�/o�ؿϷ"�]��S��]]n�-҃.�/�&om%�\*e����
�vQ�\i,|���[_)�������Ic��wCqq���V��ؿqID�(p�T'	e��4����b�����Y�qyۄ~���W�ZPQ����L��ǚk!��?��3"�"s������_V�Iyw-��S=��6�^�!y6T~���8�c8 ���T7C&w��Ԉ
�����,#�&j�	3�j���,u[��H��=���"p����w(�"�_Ϋ�"31�⪦�a�;�{Z"oYs�{����"2`H����Z��I��(b��
��8����/�}�; �tH�5�IYҶ����:�3��:
� ����h<��umLF�L�){�	�\�Co�5%#_�$��;Q�j�Wi��_�~.�|�(H�;�M%� P[�.b����=�0�/]���AfF�+;b@�Y����0 @�崥�ߴa}��i��k>ޛ��)�����'g��05�$�q�3� g>K�5��6�(eM�4p�	M�2N���k�T��>��lP��D��s��D꺱�	FK�k)�3fۍ�kؐ��`��`�	/y�-�oqѻ�QA����!�?�ք�*�6��(π���s��H�Ԃ>3��N���3fUT����-+>7��J%6�
��ɕ�	�-��9�����+����q�t���d�K��s��Z		����E9
�s���^��6!1�a�>��]�G�����K3�Tf�ݨ�}IY~<ꫴe�=��Y�������a]��I(_Z��oш��O�N[��-ukWL=��}����V�YzM>X���gz��s��籓���ܟ���Y­�3z�!C-�*�5ȱ/���E�7��`��T���)<(�.�mT�@�մ\���
!$/<��a�K�w���Cũ����Ǯ�s�G������0�Ɛ��?69�w(m�}�S�Gs��QSbV��	��9�r�眩�%�T�FZX���Y��(����������"�Q7Dy������a��{:*̏ҤХ�1���N�OFǲ���`ӒcIl�	���*\��
H�a��@y��ZubsIĿr���&�+#ۀ��"�~IA�K���Z
���rᵱ+~ҕ7����k�_Je�#m!���[�;]�������Ĝ}���b�2MC0�D��>�O���\xo�Өud��/[��6��!x�6<�"����gh���?�h?��Rp��n�7C�)��G�&�B�_�R��wF]�{�vʘi$~� �e��n	GYu�8����U.R�ϳ���x&g���]�Ǖ����|\k���s����-��>�Z����3<AǷMg{Ӟ�j�6.*VN7�K���'��������߾�^�������!'g3z��*�Y("|Wn�i�N��5��ۃ�q�$����ѣeo�7���X�$��*��a�6����Ĳ�<������l�{K�B�r U�����Pt?7��sk��Lk�f��2Ì%�ǝR��-������C� Bb���Um��f��s+�I����k��z�5�f6YP�k`$Őo�>E&�WG3@����Z��>��m{1��`*o-�B�eʗPK�֬�����nuLX��r�><�q��L$/ۂ'��ʈ�T�wh���_�X��
>U�/K?�Kʹxr���r;�"CRXdsZE�^o�"c�K��O�k"�y�2��N�(���KN���@���S�_�]��W���hK�B������/��%즐P�C@#5T,�@'��둑s�Aʧ�~��ղh����ݟdc7��m.^�-=OU.�V�⢹����X4N��	]�.Z��������Y������Eh� � ��Ao5��׆O�c�lu�t������I_z
83��E�LO]h��a�^LA΂���l��[c]�VØ����Ǜ��iҳ�ᴁN�_��:L���^=����?�z�%��;�}eP��ط$�&�5�d5C�$])��z��&?@Fഓ��8��-��M�f.$�"�������D[�ѯ�7��?)�d��+�������W�4���jc2��D�n�&�,ņ*�P��&������>��S���o+}��w��.��d������@��j1��H���II1��;&��HT�$,�Gb�8��!��V܎Ad��m�N��+�[IP����� �Z�:KGLa�@&�P�[H%S7�:Ay���]���43S���"�<3&������� "�Gγ��+S �2+/weA��`4 �6��q<I���7�w��|k�\��w9"b���X�+��`�ѿg}6�)���h���=OuQ�F� n%0����w6E�Y�l��z`��	�t�4��L���,z�հ2�

Go���&�H�뾲ɞ@�	J6�oC�:��%t:��\]'#�+z�agH b�n5f�� ��a�A��5��t�<7�E�tӭ��5�����;,�[b1�oB,��O0HD䄂�5�BQu�^|3L4	�߁�� �y�_�ᛓ�3��G���n!`ӠVM�AvF������sW��}ɘG9�|C$W5y��se�@�����[@na9�
*����.+
{�h@�|wma):�m��J���?=��ױt�ȹ�r�3��Tc��U�2��~�w��N^Xn�09��"��H8��IH�;���'���HM���Q�}]�RM�rf��i���j\p_�A�S���o�׷�uG����,$5Uv��OI^7��ezۼ��H����iLH�KWR��@��� ~�mj�g;-��'��p�Ǟ?����L���;�Ms�F>����
|��K�e-��v�f��e��%�ԡ�Gb-�Y9��3U$c	X�W'6p�N�?�oBD�C.o��T^<�������#��֭��n,^�\Ǎp54w&E2�a��	�G�!^�&�s�<*�ev���b��F٦Z8�:��Z������A����c>ĦJ��F�m����鉃��60N	�@[�@�ɑHQ����#=���M
��:U#����W��%F�70
:�K(e���(Z���8ʍb8�/��`¶>_��Z�9)��Mt��ߌ��; ���E�)�b���Jm�/�H���]o���{kgM^��w���Q�,�R���b��*`�c���u�`(�43��i7|62������-hw�8�~6�X��݆ӈ�)����9�J�4��o��"��ꦚ��[��!��%8V㈼����K�T����
GE��*Owg�����(5g���Z(}Ҁ"_��'f4�ܠ���Y��l�̭�����|w��~�G��Kf�j
�cxW]a�)?�����Q��aVNp��8(o�)Ű#��gX��S�\Zjr�� ��N�'�q����P��J���F�����|K��&�����g�C[S��������Jv�\�0P��q�"��a׊���;r��E��
��D/�8ԯ�tX��b�2��N��\YVo]�\3�ڳO����g�0���W{H͙0�$�ZMʔ����ZbPu9��rj�;���v��f�L�l&5IZ��H�2��AP^{MTGu"��֩#��zC��dk��7�[�M����'6�X�G<�!�� ȟ�� =h�t�?m�~ȯY{�ۣV��t7�hajQ� nV�-h����O���r>&Ag]|%�M�@��t�-�ܖ"���n��L�F�������p�sMD�:��h[g�oڪ&C��G��*��\0}&��G�E@�	����Ü��$�j��(��:92���3ur�&���'9V�*�9Q��}֫]�^I煃cp��
�uԜ�� N��
v�/&�&��D�c�AFBI�&�K@�~�]Ϙ$��G�
�ْ���4
Y��b6�3���PXV��؀^_l��y�!�:�ٜ9Gs��q�)E�r�2��P�Ɖ�·�4[ZWh�F9�i�BX�J��z�B�%@%w��W'^p 2����ыC�0B��"!c>KCv�(f���े�M����Kv]7S���uNoԵ�:��%I��g��&����X]c%���WE��B�K.1d�@M]A��qVD�u�nc�3��y���H�H��Ct.�}��m��Ԕ�==��G�sp�Jp>`2<a�=�v�ą�^�\�c�Ǿ7��ꯎ�&�a��>���Hjm[�W�l��s _�GB�H�S��3`||?:��t�`�G�}�(f��Ms�$yR��՚0��;�?�T�a��]���������K`��C�����1U�YSW2O5Њ�����ܠx_]�v�O@�Z,�i^�����l�ԗ���B���Lƛ����6�'_S���!�Ή�`N�u�ɥ�j�������9�t �zk#m֗�jeڦ�F�Mb���h�!������{%v3vz��ɩ�7�w�F���CCc��-��o��\_&���W�������-@z���`/����n��"���;Đs�ch������'
��8�F!e�q�?��xЖj�w{ՁN0����j�E�� ��b�?�?b=n�>~�W�9�L��cRˎ��ڒ���p����Ъ���Dљ�0��z�z >��ƞ�&�U�`���]�ij^-#��9�~�2#�
v���R�"�t��h!a9�N_���&O<dP��"{a���7��e��G7(���mN�E|B��"VO1J�!�=��*��+��G���l�B����AK]q��2��-Ict�$e'�^>���+���Ӝ1�X}���&�u5�͝ݻ9k����SX���j��Z�2y�AY���	��B ����B	��W0O��yp���(�bwV�=�ZG�?�����q��<�e�B�9�v��B1ٶA'�Is��Z�b���SI��g/Uv���Y�k�aW��Ny��eXn�`��e’�����R�v/P=�~S�g�9E��SM>�FZ����i���w����e��qR�����*����E��0��K����=p�{�mwT����wB�JfX
�[���z���+u�s�w��,��B.��!��
�u71d,zŃ	��,���$+`���鬶B�D�U�:���3���ȸm3( Ӥ�8'�@��K�y5�u��Ϗ�KCD-���P�=��� -�pL���;Z��l��jȼp�����~����s���m�\7��Kr�PB<�]���>M�1.|��Cd����o�K�"4 W��Q �$<l�:�cH�~b�Y�Z�T)��S���0��\��>�.��y9M�̓�Mߩ����"bJըs#i�B��x�M�J�[���E��$�sr�F6H��J�����t�����,Sv��#�]�n�^e�A���D^$�a�?%�/{�d}(6DL2,��[��=�><w4	E�۝L� �����g�`�P=�o�$(:ƣ��,CΞ曝*ѧ�J��`z�B.�.�{A�}^��m'�C�|vg�s�o��.�iT6}yq8 /E���#�j���)���q��\4����b��<3M��H��A\GM���ԩ���l��y*p!�Vh? �{-�-�0Z�u�\������N�����T�RxV����]��2<�,�D$�+b�d;��_4t���+J�|�v����]#�D�:�,G����M�?7��+��� � �yOU0P�M_�<�8��{�0Ei�7bЭR������i���=�NG�2�k��Q�[Җ���_"{�����1�&�������z���`�?zTb�Ѯ�"O��.X����OW�j_�j�4�W���Hb. �K��Alj\�m�!���D�a��VB*D� o8N��+��HhlWyH�8��h�w����kA��)0æ�6�@l�����Im�AcG�E��$D'V��=����$�81��2w��������?�д����(ʘ������ gdw���������0Aj���-���aD�W�K}�@���߅|+'/��9"�S���?�������\��f���5f�Hlrג �*�h���d���BO�K�ZE�����9��Kx��bC���!����~���Φ���}��KT�J&�)�W������R��wV��R-FD����֢��[Y
�G�%���D�a����*mʯB����%�AJ���,����{(�$
3A.���ʹ�0o�a��J��T�
�L��4�j��\_�����1q�y�"�H��wt�4�ܹ!�t�&�;B=Fo�-0e8,'{�2X�|��w���[�P�Xczi�P�L;&0BӇtf6q$��<мam�Щ��5
:�ⱟ,m�?;j�xZ�4"�]唰/�Q�����|��������Ҁ�L��a`x��z�b�E�|���� %�m���M�B��
#S5�c���)��E_4&"�~�2a<i�����V�ki�s�޾��L�������<��^I��7�H=�a������܉Z$7�׳��	kz�P �S0{\L(0���2��I*�p�?e\xM�0��倪i�H�V���0c0;�S_��Y�M4��Eҽ�C>n�����YB�wt#k���2��kz�%}�P?(dY�u� �8� ��o'#��2O�c#�l�Ϙ<8�%��Q���Z^U��dZ(2�t(�7���ks-�@؂�S��!4YǜT�%�{����a$��H�����#)���rvlA0m@�KU�����Y��,��ԁi�g�T�MZ�? �������LQ�{�|�ZEyp9ߞ���7�]���ȖI86l�Q�;��g��n�������#;�C4Y�PS�$V�	��K�
��:������nI�@&�E��x;�*i\��)����0w�\18�=�%�_�B��=f�'��u�S51�{�gS`����S�R���˚�N�;�������:��"�\�f��H��s[<r���Vٛ�2�#.4�ͷ'�З�옋��U/sO�N���A#�[r��=�RKjp�zR��>(I/���-�'�"�f�J�����;�W�Os�LR���ä���y�����1`���EI���*�[��|ɞ��C�o衠g��
	���(�'��qzY�"��%/��$�lp'| 9��ǶN\���djJbT|�Jt��B�tkɠ�ru`Y�g��sCG�4�#(拦:%��8�����.7����$�6z��:�Aa��$��.P�Y=��|E�Xu~v����1�B���U��C��Ж�kɊ��G���$6�h��+^�t��X�,��@6at�Y�L�l[�w��u���R�M��pB屙MҾ%hS�  �^�G��{�A8�>@��O솤��<(y�Ш.���)�S���?y�m�q���+�δor��K6�*J��k���ҒB��c޲Me�~/���x\�8E=�uc�tW{�7*��"�7��V��}u���#)�9e�p?�WvNS�N7rMT�Pԋ3OX�Kr��F�����v�@�����v��}�F��{K��͆�Pӱ<��"N��wq��.Md=��$@��'M@�
6�����c2˝z#!�� ]B7�!Ep���sۉ�zG"����o��R�:�@��N��#�@'%/�;��L����c]��J!��;VW�e����}�Skktz[?# �ܪ��>���&+0�~C��z��z�=�X;8��6�4�'O�%̏�n�-�����\���ľ/���OPTs:���x<+Ks�i1ϕ3�
��gd��'xRF:^�e���Q�U�_�(
�-��wo�2�X�95� ����C��DH҈���={j������@q5-��c��.]�fn
��	��d��.� x�|�U�sM����~vW�ɖl���ɻ�7 ��%�sp����t�O��O�b�h�3�ƃ̌�y��m~V���4�p��Zm�9���?�$��7^���X3�.�|�?c89ggZ����YU�y�3���mDJ�&���R���-c�F���Z���)�@����%��ˣ L�iv�g�Hj���UӉ�Z�^�R��[����ι�Hݭs��+Q�X�����}���W�5�!F[�����y?������|5����x۞����2f|��u��I�}����Y�`�ḽ h��A�I�����>3���^v� �w�D�}�Vz��Wcl+�G"����L����ː���@̟�b�6mh�?�!c��Z,���y�Gd��µF杦D�̳?��n2��l�*�Oz~�=��2�4�&�����=Y_��S�SU'��29F{%�B����)��%����A�>;V�T����Є�Sq�<�{2U�!@\�f��������p�g��AD;ε@�X�LPg�ȫ���c{U�E��P�A2.=SN<Q��$A,e����w�]�uu�9�<Z�z_"g���ۜ��O�Z��Qs��!e�^�9xϸSG���K��y̴7�
�,��Wi��g>_��q�k,��G�ߡ�ŕTFF;ɦ����7���(�g������ep�T��g��������g�f'CI�\)����x��^�9etp)����hR�������|�YGk��3F渁L��b�!@�,j���������IvZ�9��~̘�[p]b��	&x�{D.�x�K44$��·S�R�f�����cd�[	���XGAS:M�s��q`ҹeC��<�Nx5�כ,q��qӂz/���a����L�1�C8���a?�_�s�
,�$9��Dyl���e��|]'��)A�$4���[���
�M\�s�����\�>1��i}cS���i)e�m��D0�a� ��.B2a;���hj��j7�1��������F��NZ��U��Х�7v��C~w�J]g@ߵ�M�%��D���K=�v�v�ߡ ��B��V��lw��7|y�x�����{����r�B�G�y�-+�����*�D�iP=H�/(Q㧅U�a��?M���ϮC|�����&u��1�goK56���3�?��|5�ӄ����xwc�0�.us��r�Ê#br.h�Y
�\��8ޘ2�gS�����en�r�����T)��T���+�0��X��QW`@�^�S��r�l��Ⱥ���-�Y�l�[r�˷���e_�KCeB�b�P�H/T��D=�I��� f/N:��CC���-w#���Lf�zh,�� �e���pN���2)3&pGUtWW|O��h비���p=�/`��e�*0��(�ȱ}�R�J�mf F�
ծ��)&�i2p6�K2ՈQC(�y���@����1P(�z��5��i��&�{�#���HՀ$=B����(Nxm�Џ{�Y�/h�Wl���3d �������*��ꯃ��j͓�j?*d��jhg!�c�:Ɓj����ܙ߄�[-h����K������8e��]'���o��p�Yk ��wT^�Qt�4zlA�'�שW��S]w�-�wN���b��x~~@��<���@�^��n����t��O�iX����{����~��n찒�w�=島V&n��o�����.�g
�ɛW��b-�O��r
�Yꌰh�$G��E`�@���/J��b7 *�����!�F��rL����K"�2TL�?ۤx�`��ߴ�u���Z��ߞ2��+��Rs&$w#��X��B�5�F��'M����,h����Wo���FU�]��glDu��RN�J����l�R�b�-�	�0O��9�4l���4����,))tVc���n����ѳ���>�M�#��M�с�$�|7W�P����kGZ�~�~In����|{N{)Q^��λwA�VzR���Q� 	�erM"�Ϸ���	/P�=t�(�K�'l�{5��b���N�^�q��~�V;07�-��ė��BG2p��f�/+e�~�CAk}n��AvXAl�������vQ�K���.��� Ck-�5�Q�G� ���5��g�#$ض���r��5�1�<���]��,�6�*è7,|V��?ٺ�>���<l9+r�=o�F����"$
�[ԕ&�����kc.��ы����4h��x�z ��~;o��^��=��'�V38�_�ʿ϶0�1xd����禷#���
>:����3N���`���ђ��/�������R�C�q"���w�t�#���6�$��nDxc���)()����m��S=�zGd�k��fw~���+0T9�$�e+���p�Wq�Z��t�ő�a����`@��WD���b�U�4N�4ȅ��X�\ǨP	Pl0M\L��~&�b�=W�T���$`�s�7z�э���A�k�'�D��-� T���5���~qɕXsA/%��!���5�Ry�h�S�ˣp��=��)mO�mV?��î�p+��`,���l��_h)����tJb®|�8Bע��X�z�m�QJ�*���0��k��G��ی_9��1����g�����*֩�����6l�q#n���"Cf+�7��>ע�S����5�_�5�tE�wo�P��#� ق��up^(��xy1u�yw(o,E�����z�bB8hC���������ԧx �!e{)�O��������� {sl3�y�;w�c���[x��k���+����>���2� �ljMі�m$�؄(ͥ?��7��`5�92�٪ٓ��X�#[yB��� ~<e߀�����`'=�(�H�I����<�`sͲf��"Mb�J�M��I�:�³�2��)8W�*���9�
|=:g�=�^`1*7{_��*.ʝ�S1����;��jY�J�e��~��m�3ծ���l��U4-U��������k�/�$����
�LCsJ���F�%C���2n����uc�a��͆!���)�szU�kW�[���S+�Hr%�;=���[F�;-�q�m�5���T�}�4�^�e��멺S��ԭc����8�"|d��e����)���+�Օ:�p�z�h�QVl�=k��?<�Z�7$Z�9���դ��$���u�V�?p����'�]xcd��·�t��.�������Q�5ԝ�im"ij���ہ\X@�x�����l��?�oV��b{l���i�LK�H�,Zv=I�S�ӥ���DE����4;;��?����lQ��Vk�D���"�����E���cA�MU2��C�s
J#�{$�xl��F�����)�sl_�+�("�ew~F�%np[��3�p�Чb*W�I(�V'��p�Dm��jY ��;�W���CG�X�'��-Ŏ{�O��_υ�?q�C[FY��8ʔ�dm ȣ�d�=�|<4ufgW��	A"��ur��o66́����&���>��ߌ0p�����3샃,' vi��N;1�kbo�i��9���/d3��S{�XQ ��YMG�<��GL��߾�D�µ؞ЍZ,*)�z���Q����s<��y17���΍��<�^l�vQ�3�l������XMuF���8��6<S���L޻�:ځ��'��.����n9�Z iǲ�X^�ڀxg��Q���18�G�[����$R�D�W�� j*>.uC��|@d��͚L�ߢ��vAy�q증Q�A	��R���C�N�Mi;�]���%����)}AǎJVT�@N��
���Z~@Q�k�x�'Œ��q�'^��FY:�A 4�=7�nOfՕ���#}��_o��X�v�:����T�i&������T��IKZ��&�(O\~��	�k�{%�N
	.��ҢE�w����� |Y�;�S�{�o �R���ݺ��'W��@[�����7�c��ea�!��WΰXX��u@EUA^P�K��sW��5�e��4g��_��"����7���s�h��/�G��1��<W�f&2�?��r/E���>�2=Ӕ���t���(/�%��m�n=�{� �i%�b�ő9?��rcn秏��?�c!�fh�j�UZ�
T�3����˂F�V�ȋҔe{�;��l�>!c���{v9)eh]�#\sb�å���5:�g��������"h-��9 8m9[׬)�$�j0�4�8E��0��3�I���%K�2E�*O�,��������K�,��Xs��BL�0�t�����͉\u�ث�%��4��+�L�󉿙wmIFP�f�E���:3p�PFW���VƐ�K=�:�j(J����u����\	��-,
8��A0*�,��SJ�MWI~��XB�]�]�f��k�*��gr�Co�{hE�-iKi�d���?�^k5�@�U��*�t�KeO�r;('��t�S�҂�?^!��$
�<0�������+��� �.�׸��}+�A訠�
z��&�=���&�-��K]���_]j�C�4޳��a��#��N��������Oޡ�'(4��G[�gY�׍��^p5���BM��y�߄	#��C�/&�;�����,r��݁��2o��^ϒ+�"��R��)���K�%�#�_?5)ֱt#��p�����Ld����I��q[��㡐y퉉D牏�@؈*+�䎥�3|��:@�3��������X
��߮�?ٕ�ݮC��3R���>�ܝ퍿p3[���~��Mb��[��	�H�iʂ��3���И#����z�e�|mP�^{� ��W0k��S�7���6<��߆��e�����J_��GGox[-�ҏfcYhU
;d �Q��gg�w���I��ꑨ<���|'�~V`�V*[8�+�뉁N)��N>�Y�H�M�1C�T��	�E�T��@���G�ß�A�Ew��]RN��^ʨ�y��K���W��c;��7j4�qNSM�$�<�G��	m���?;�͕�pZ��h^M��]-tZ.(���/�B��Jdnx������ �h������Ma����.�p��(�C�T�'G�y �=���[N�ić\4 ?���Ӫӟ�ԻH9<`����#�x���S{���dy2T|ݥ}�^����}vT�ȬzZN9����Ƞo|���X���3HTv�+�z�b�k�n$�5���]��U�`Q��u�n�ô�c,��v	����l`}.� ��+e2��H�PŶ.���~�/�5f/�.
K��O�wM��1%���y�p�iIi5]2� ��FV�B2<3s�V��3vv��4���[T�ƗUtm+�WI)A�Nt�R.���s�5����F5���̐ʓ#�vNe�g���uO{�Lgk>��I�y��셱F�v2��G/�4wk��0عU�E�pڽ�O�Nt�O�H��#�$Av�VǨ�'�H�@�J+�{N�E��V��3�AbL_`]ZX�y�,�Xԧ��O���@�@3fH��k~+�F���n���ۯ�A��v��@���d�����f��d�Z�g���lX�b�#�eP)(.����ٕA�Up׬�Z�|�қ��+��F� 	g�'����]mȤ�_�[�M����yhK��
a�S��n�ڮ75��"]��](��;�5
80�_w�&�y����N7;,�d��a~�-�����F�mvy�QՎ�gCr�Q(���ۿ�i(��O��E��|���,H�W��Hά5��Mb���L�����6���?�:���U��]_���ۖ�&�`�Wr�����r�^w�� @�����;����m�9C�!|��Y���[�F�%��S�'��y|@�������֟B*w�P�&����C^2���>9o����:ȍ�9�ݪ]$Tu�(bI��!��ʨ�K �2$!����Ӄ_�S��O6(�|I�����֏c�9k��v"��W����ZP�J�^�܆�1���ǽ�d� 6�a�	��i���������$�������.�P���2I�?��J���=�u�XR�C��Y�k�渦�v�F�$]=E��;lu|4�?UEn��W�9�*cͮ��Q���%��O�O���y�ˣpI�X	���Ӈ�bH��Ǔ���,��'B(5����=W��3%9.�׵2�|�H��[,;
J�S0��oQ���bO��h�9=s�-"9 � �������`Z��\u���cʾ�4w�,�e·Q$]J����zE�I���`�D�!h)#��y68����v⛲�Bq�hwnJ7g�����z@���W��2���m�2p�?v׌�j<:Jb�6w}*��?-�`{d���5Q}g�($�<.l��� ��n�w0��EL��rc�g�*�j�:U�,|U\mK��N���򾓮����ٔ������Wd���G6�h�>���xL7>l�䯣��������9���kiז��%����T�x��.[!�{u�K�U��H���OlfIu� .)���(1l�n��c����غ6ڛ�4@�>�#b����(b��6�I���d �����oRȴ0N[ke9�Ex=��O�=���+��?A�up��r���o�m�`!��@�4���Q�;�F�������KY�Ω��?=i�0�k���3��ʩkv/�H^��Sm�;苾.��A��;YhX��o��,�ۢ��su�u�l�Q7Q���C6?�b��^6r���z�1���(�fFF���29�!E��,}�ǙV&���,��f�U�^�o"E�5,�W�b�gS����So8:���u�?�������0Q<Ә������ã�p��f$e�E'�z�����)���ߒv#�����5�|�S��0�����-�>��tz^����q�/&#t�a�<DD~&�]r�x.�R����3z�ƶOU���u������M�d&�B��V��Oˠ�����x�<���f���z[O]�iT@ƺA��_J���@hi���q�n���t�C�b5fv��ƚ�����¶��`�1����\vV���e�c�[��kOo�v/Eɦ����4�('�hM��<��X;F�Z ���cds����O��	�{èK��
lV����Y|� ԣ ��=�v��vd������ia����fb�Yػ�?�N3���i^spS�1ASx����N	t
zFɒ?1��f=��A.N��t��:���a����\���Bbb�C,�T㆜�:�%r�~��x��^䟲���[�	����}�no��ҩ]h��⿇��Č�x�F?]CX��ޝfy�AN�=�_���pl� z��4�v�=F4��"nzX�7���%��K���.��gA�g�v�efbY0��{���]1�16��驗I�y��1�V�%E��߮��zKбq>;�HҗF�J)�m1�ɛe|~&����XP$������@ap��a�k���L�J�vZ��c��(/��������-?�����%������߇��~}z�ƫ�k�E)"��|��o:����8��m��9b���i蚑��2��>�o�a�+��^�/3W�����-�Nh���5�� {ɇ"���h���Z����k�����(J�qV����ۀl����wFoʂ-��@ö+4�\����#ܝ��������<��^�P�C��Ր}�M�w�l�i�L�A
=��c��m#�,;��g���2�Ӹh-�(�jg���Qo�D���*��'��������>ϿV �yQ�����	c{}<g$�����l�����e;$=,�:<��8Ҳ��-��$�	'����B0:����D�j��'����J5��3�;�(ni\�b���+lDx�d�}�ir=����دY�S� �q����N��w� )����OI����+����U�ʨhi����,��R�g���ɰ��d�Z������H>�YƱ��ؤ��,��F�E��5l��}���*E�9Eɼ�p�5��fzQAM�����z�����0�2;�`//�����hQo�y	I-�z۱
�����H���{��ߝ�z�)7���@F+~'1*d�I�+ �[ɳ��+W�O��RZR�,1�*���Q-m=�ɾ�����&���T^�yQ�dά.k��@��^��z�I�f��"�݅�"�ʶ�����C�݇J_w����[��S�A��oPR����o�s������CJ1�����| '-�8T!��Rf =���Q@��KmE٬�	��sЯq'a<N`��)��Դ1�|%�G	e��F��ᤥPT�j�2]�F��WG�h*��������-�Ԧ ş�1k��w�����y@�=JX�P_2�k����� @1}��5���1.IG|�69�>8S�N����x6��0�h��N�PDl;�b1
�:�����������I�a���ey��9�ݭY�J�3�_P���9��J�F���GԖ�đ����ѭ�b��%N���ZWM��� �����.2#ӯ\���0D��C�1����P�jW@C���l'v�6>C�=�%#��R��PQٙ�V�Ԙ@��G�JH�(" ���|� u^���nJ��,-k�t/
~�
�HP�U.�B�J�_.T0�f�.���s�x)�H�1Ga$�=��IN)*�97ú���!И�����䖳]�Y��E��gk����ЃR�`l)�ؒR���E�U1$�˪YA�	�s��Bb����Ů�t=�O��`�Z* �o��º�e�v,�h���*3bl*K�!�2E'�����΂���o~�Z~i�����������j��'��gs�V��\�L�Sө��F_�2!�ܝ���+��nb8[���G�
�̭��|ǹ��X���pUP�YD;ć)�J�.��4ԑ�kZ?�����|��ݴ����RM]g�����r�>۞�qI~��祺)�md�2�`O����?:�f�?�.��S��t&�G��G�~�s4!����Z�����dF;�e�M)�'��US�(��D{�	ʒh��AT��`����=�{��|ω^$O�m�����ǜ�-�ޞ�l���о�+f#�[i�<���#��tM��nC�� >Š��V��6��?,�˃4��EY���2�W��g$���J�4*��:��U#�˖(��4$�2��"����礗L�5&�����5D0�5�cUA���f���Z~�\NUi*=�V�46�����)#�z���O�*��+�S�j��QMֻ�<b\���9�c���B;���������v���yh��Td��ZDE�ǒ�v�>,ۘ����� [�w�����G�S���"yj));�+1?F󡭘Pv֐���vw ��
�C����.��oP�I�r(��i����:��C䚰<�]~�̰\�a㈮�맘��x8�R/{jayj4�ab� V������ � � TD�{CJ�Ȇ�)��'��y�\=�[	u/�.����h�PCz��6;�a�r�+������J��XPE&V�� S�{����+y�Fj���^�S�#���[��\��"w� �"=!q���|�M�g����U!��둝�V��O��M�H6� �Y*�2�����'���G9�y�eW#��g�l8F�xR74�&%-����4����n��Y�����Wl�lo���*3�a�YGn +tHmv��9�(�I� �y�
G)���6x ����������єDLl�]��z���
g�'r0�J^Ƴ>�4�E�O���>�OH?������!��;��DE��=(*��]�/�b6v��-����(�琙Le�(:@I�IWC��OW�z����Ԁߑ�c�DIwB'~�z�T��{?l��ܺ��=]q~�8�*6|�n�Y�k��|+���cB�k&'8����������p����=��(�-�@'��'4:ҟ�[.��E�.q(�]���Wd,��.w��`<����r��m G�d�7�c��̩�������⧦��B�Y��K��!ׄ�<��(�y��P�G�G6h��O���	͔O[k�၏&�{�wD>-���Jwv�k	֓b��߲r����Hqf����g0��f }���NF�������@��S%�� խ=�U����@>��S �dT/��M-�n�2G3�GIx��H��X���H�A�]v�k��Ǩp�e|�^��%��/��Đ�yM�Zq�7#D�*�Fz!���ʚG$kE��X�t�֍2���/���l�*��uk8�";�����}6�C{�*gV�oo{�J\>KL<ťĄŬ�3���= `U7�������c�Lk�yI O��8�������`Zu�j���l��񯁉\۳�
J������bQϩEP�AL��m0���Z��V3��̓�
ҵ�ˌ�D�<5	.ց�����y<`���C�l���Zlu�U�*o��= 
ޝ�\�Jn6�pF?�W���$�Q�-]����v��k�4M���( L!�e1��C?\/�ÖW���Ğ^���R�5_��y�q�d���0��'9���{9��Ésd��')�	k�Cmϋ��4�jU8*�o�I�0�\5m�+��~�� �ǮV�CO�'���2Z�6�?F9�ʱM��/ |k�A y,��Z�~���՟a&����������<T}Dk8o�]8��)��l"׾����+�'�L�n�g�d�|��C�
a��l�K���}�wo�d� >�����W�����b��]����@J$6�Dnm0�9�<Rʯ`t�Ď7��[�|N�*8�?�7n`jE��e�J�l�x���W�b7d�.�#��ݚ�p�)��(a(�(pb�-.5�^i�u-XC�ڋ!$}�OI��� ��%��<F���8��)�52���7րK2�!3Gi�4��� ��*�;*H�vɝ��\����_�1�~ʈׂ%�-��ބ<�����]��c�=�3ڂ�L5� |u��Wo��>M�]���aƴ�q�e���Y�'�"��oN;�f �;��U�[�δ>��lI�v82�����@����Si�ך�c<�eH�� �H���ޤD��b�E��)��~e�*�Z�e�g@.U��:��7�鿈��D g�9
�@y�b+3��Њ�#���o�^�c��e���@����}\�9(w&�B���+�������W�%���~u�4W�b`������p�W���Q԰���P��-�J/���R;!��i�n/����K�[7��7�
t�f�x����yڄ�J�$�pN�}��A��Y+��T��O�x�s0��p'f/��_�M���[�1氦���A ���Pd%�"Ct�Т
���7#������UH�rGrРe�Z%�Wo�﩮c�N�ָ���2�o�g0rx��</�Cx��0gZz�� �^�l���h~~&�m����X3rH)??-��_�;o�G9ʯ��՜�������Q�����w�I57=��q��c5�c�8��<���{'jN*d�8.g�,�C.���\����ו�d� ���C��D�j,�"��=����d% G �%S,���3������P�UIK�
2�:�V�֟ѢB�{�rn��؞ȳ_$W���C�|��m�XB�k�Jgp�zX@1�C����m.�1� f� �5̷=+��V.�\^q��&�A��,�J#�]k�`�d����ϑ��I0�I�����C���yx�ś*���
�-v��u��#������V#_Q�}�#̫��v�!�i�È"(�A�o>:bQ��0��rV����I ��^6)�;0�g��#�ߪM������˴�ʀ���4��y�X�,��<T��sj�{)���uс�Dѓ�*LR���%
�3���X�����2��5����0����K�$ׯ�a�D,ƶ��AϞ���h"�k��Ť̶H�����l�+u	��J�6�7�~�o�j23=
��F�Ȋ*�u(��C��<S�y�Z��Z���)#T�J�s��腑�ʡ���~�$�"�l��x\0�F��%Us��g�l&���t�c�ѡVK[��R��G�Y���*s�4l��6�kn�H[�u�p�ގ���q;�Ѝ��ع%À�6���f�,q#>I�B�ܡ漹�B�8����P:�3����6��`��b�ӕ�a��+�-[�n�N���L�~��~m��T�8p�(��f� �&�������w�M:��5��n�\�S<*/s��j�.�x�A�_Z]��v�5`<�KJx����lp��"=g_�O$�'���4���C�����n:0]�ڃUą��-�#��4��U#[�f�"8f �\!���Ț'����[%깼��/	���Ju�.�/�F��g���R����.�H!��kl,�qwDK'o�)��7x�ه�K�n�/�?<�5�<��8������a�[�uuSv����<�VD���.AW�l�DZ�I���GW����.�n~��^��җn��B����܈�[�ڱH��.���`:�Ms0����4<,��ӄ��Y�0��ԟn@_���x����}��S|\�sН�����T6/w�9��Ǚ���2G��3�&:�#�%�\4�oq�_��#��LKV۞Ԑ�,
N��MND�9��;�oN��Q,6��w�bW0��k���md~[~a�֜M�zn^�$�@D+��< �t��W�;�� ,&���o�V��R��wX(�*��|�2�[-��~i��akqw�Ha�vi�u�M<~Ҭj"��(8<�@fvbǮCq��i�,R���ba��=4k"�>�by��E�qx�2��{Yw5i��=�)2e*gW�=�Re�30�C���};�V�
w�I�o��J�0��w��=��×T�"���6]?n���Hg���2�7���1�)��M�c�֕Q��Dh�+2n"�6M��.�((��Yd��_������IiR���.fSo���4?V��ܿ��^v��]˂�	<��K��|�:%b���i�Ñ�3�Q2�0Jz%k��x��9%P~��e%-Y}o`�~�o���x�Y��1c\��w;$����cH��?e��r�W|t,�l��m�OZn'@��
�u,u�ܴ�r��kg����T�;uL����*z߫f��Y1��.��N��]����u��������|<M�V��'�0�=H@��hSm{j�?�̆@�w6m�����j���R�*	�RضtW�Vig5��k3mF��Y��9d�������3������o[]i������t9^����O��E�g��7�Ui��T>ی�z�)����߇�[�`'�)Ɠ��t����,@�j�X�Qr����=�4?w�iu*?9R\O�B����c&���n��L�x�ˮ������r�;Wg*�C��v���Y�"	��Cj�j�f�����#}���l�T�ͦI�v4�B�������0|��8���cq gi��Ҫ�6�fkG8�`;�
�f�<�
��6�ݎ�Q]jב<�r�:[�v���b0y��������G,��k�s�JVƤ�b�iY4T�3��ue������?�@�C�0�Qc$eÆ�ɜ,槾Eʏ*D)��3��o�ªM2=�Q��B�DiOILs��ǾY8R��,�P�D��0C��\�M�|��r���Y>�݄��x�i?�K
�]�P�pa �n�#VhLb��V>�T�,��2�B�bLB�~l3#8�j􉢰ύ0e0ن�6Z*�M�Fk��t���ӂ9���+X���9d��$��wyx�f���h�|
���:���<=e]^�-���kE��'�����cK5�S@�r˴��k�q���%�iu ��/�Ri9�������g�p�٥��ne��ɪ.MG�/��S ~@�tn�J�/�.��s����匐x#��H��<��.f i�*��l�P+.E\�����E��d��#���H�|4>�;�r,�h��&'ݺ��������~df�Q�B�S��T���g�gid	i�w���^�����`�U0�St�_��G�-x�c�T��t���gU�������#M	�����?ʆ�����dt��� |5Lx!�m�Q$�i/iO��Z��dLB������Q:��fP�{E4%��&?�P�pV%��k8�����֝ �W𐩌,E����$ك�Ȏ�}��i+��A�������g�־T����38��o����o���l�F��|.J�<	�-�'���#��.�B���|�_�	��/�|w;�<U�wG�����6��Y3n�B��i�̓��d��U��ɥө�{��ֵ7�߹��j�B��8;gG�t��2z/u�?�o����(�;������0����:b�����g�h5��1�O�}�����g{6[�K_�l���n���UE�)>�
mLMA�x/n�g�,*I�Aڞ�+�D��C=r�Q��*�ϔ�DE"D�_A�Hw�r��.]���ӂ0��l�l8x�!Ub��u*�3���ڜD'.�3E�R=m���I|w��y*ٞ����N�Io��N<���>%<bҁ���0�Bk:�@~�|�
f����/ V/��V���^��o!i�%V��˒2D�r԰�[ř�5Ԕ�W��W.�LC��]���F)��(�~���>�A�Fn{���� �+��K�zI-�2ݪ����Q4	�m=��gA��'�>�,֚�I�-zo(��?��=�ˎ����fk>��9�<�z��G��3ws���--���0��d�	���,��o���t���P4���Dg�S>JQ]��XE��z����GX�ȓ���y*lu�Y'�)�T>�qg}�奈s�`�qM&�2,���	 ���E��ֳ=h��槰�#�g�n�ntV��9S�V�l�� _sf�t5!���A6���b�ԓ�.}tS+�=+�,��"�F#�`|$h׭�v(�}Dr+ �p�)���ȼ^�h�#q�\���*E(�Z�}�
z�L�%㟞p:���Ou�8W�8�/g\���8��F���ڦ���b������pgS3yD)^<c��&կ5V�!���i�.ؓi7u�%̉~)�@�6A,�{���&�ի:���݌o����!�'c��L,�D.����]>���H�#	�VB㻡��h��?,Mm��� 5U�oD~�1��X���7@rS]i<�#�4�7YT�*¼�2c�(5'hx�}M�E$Îh�}�1Ur��g疵B)�5��׷�S�L8
GJ�j���R������{`���1��|Chvì�x̅�$�eʁ���s�M�h��u��*K$����s	Γ�LL�H�z������eM�Ӿ�ïӤ٤z���<>E�{���G�~M{�G�#?e��&�F�*����z��2zd�g=HM�Q������29�����iB��u�qz�!I��L�߶,9Z��x��S��o��-:�"�����͑���D!��.~�Mm�5����R��"��t�����TKD�~���e"�x�a�tY���8R�<���b����ƭp̤��1:y�xO��?7�����]�����v��n� O�^����f�L?�DF�?b#�rh�K���2;9"L����IDq�3<� Ԭf���.&�!�<���'�wEz�n[`Q�q���Q�ʀ�[D��"��5�� �|	�gPy-��	e�[��x�P�o_����/�R^��3" ޭ�Q���@����g�)WT��a�߄L��"��0�e �.�^����j�6��y�ѐ�?IA�Y�E(?�,�׬�1�O̊��x�F#�M��$�����?k�(��=Xg�YA��" ��r_�~���C������P\�beX!�ED��m����']�ͻ!�+N'(����v,n� UP��ժ���P���aA?�:�e-;]���������u?�n�:�R�w��i8�B����/���'Uh��i�P��~ᐴ�4�d�[tҟϚ�lq⨦6Îx�:gb֔�T�SRT��
�i��m�˵�hw+�.�cEx+T��<�Qd�h���
���2�^�69;}��V�E���rCb��4�#��b��F� �(����݇�����	���7u7>Qъ�n��.�3`H D-�������$��>��5x*Wˌc�FU1_����7�s�v��q�K.��Q�J�fC�vӇ�!�n�Vޙ�r5'�b��Kx��=�la..�����ȋ�|�(����X���N8nc���㙊��3ݵQ'�Ł�W_�%���R�D�1���X�<a%��C���b�ݓY�w�;@��J�G��$�n_���w��ʥMQhgmOw6�E,�@�#U"ң�;<�3x�T�ܒk�M�Mfh�n*��M�)D�_wv����T0~��.�A��"��k�[����S�.H�Ä��\L�Z�5��H�.�HJN1�'�4 A��MWM<�ŕ;�)�}�2�jЉT�6����z�0�X��XD?(�XӲ_"��F7�w8��2eF�u1H2T:��G|dR���+>B����ی�ׯ���ģg������'p��_0kL~��P�k#��H���D�ŵt�����έa-i���n�2I�Y� v��Я�f���R�m��跌�f���<g�H
~xvkD�\���dak�a'�K}�L��W�|�̋y`�Ԑ\�h�ް�����=�I�V��z�(��PoMs*^�ab���is�0���n�[ ������@�t����/<A����c"�{�����JJ�=�*�aM����m�����󯺥���l��D�d�C�1U�������	��'��%���gQ����05��w��(��$p���>�a��!R"S'��o%����I��ra�C����ez!U�1ZT�_�zъ�G(�*#?@qmi|X����*ؾ���O�Z�Tل^����Qb2b����	���l��1����g���<�uî�-V�w+v����y��/'�{F�]�P��
��>�����$��[�ߝce�!#DB��w���@-żji�7/����N�\�A���?�:�֣�|n#��zН�L"�Er|��먩n��\l�]`<��J¥%
����� $7�Đs0�
Z�Uw$���jS�Z�9�f$u�y�:{B�ڂ��ZC�绩
̨xg�b�<|l�s�v";�vXS�$�L"��h�Ä
��D�hJ��|EZn�|�T�V9�g$7fh��k��|����7vy:�R��P�;��?,��4�{P�ȵ$f���{�ڸ~��F�������oh�"0�t"�2�^
h������Yn�N wr����O7@ré���i�k�vū$ߒB��֝�Eђ�fm����nk�mW��f_�U�տu;Cj��IL�24�J-b�K�l>�>�����+��Nڬ����K"�����j?��]-4Jk/�b�9�,n1���@��~�������]ef
٪�,[��9�J����u<@�z�/6���H軃/�S-s�T�9�\���!�j[�`DHf����0��%���1(��9���~7$�/��߶�'��A2o��_~�q��R�<,6���>�����Ű�®�·���M��Pߨ'd�6�:,�r-S��|/����	r�0/�[�t<ۻ0$76%��o�5v���.��S	��@*��Ȼ�"<'�0��#K|,�|
�ϬӀ��7�B���'�;��ߘ������iEqy����l�M��mS�����N���$��ccT7��h$�%��k�@C�l�Ɋ��ʇq�q9�H�K7D�3��pi�M���NJ�����܉c�*RF�<w������5Ao���� �B�Y��tR!I ��S4`漯;AZ�̔�̃9��[��n�T�p;g����^�x^?2\�h�^ӓEm��ꩾƮ�Z��g6j��~���:�����z� ���A�+; �X�3�ȧ��K��U=�5�1��A�*�[P�坢����*x�s�tƸd;GK5�Ŧ���+J�h�U-+a&�f��`��Ǡ�2�yȬlPJ���\a���h iɢ1�|����7u*�4�@A<9
p?"iV���}n�Й{;�WD�;�c�ͭ�W:9��S|+.>��B�Ȝ"�2a�G��ŏ\��p�z�_D��'�&ʟQ���dR�ɣ�奤H�j]�`"��;'���ӌw"���{�T�v��s2�V�t۲p�p���V6�q� tb��|Y7��"�6��bлww�I��i	�mJ�4eo���X�E��r%u�q�.W�!9
l+���N�fk��'�?��-��;&S~>07�\��h#AIv��,�\��9����|)xe �T^����|�_���Z����B�C�]�T=��6Lr���W#��X���g�oV�P�Bo4��Ɍ��∟L��fHJP��O��[�x�Fk�xͨ/�\�Ts����D�Jۜ�,2��S)�]``���u]b�H�;�jV	�kq�A�kn��\�;ٲ0�8\��� �mI��PK)�]�p�#�t� ���a�88ղ���DI5�M�s�#�Wz�0�W-+���Ic�2p��ƌO�Zu�{�rlygE}��~t��J'+w��Bk꽖��m�v�\ve�	���+mF�Tד��+}��^>�P�� �zi}1(��d��Kn:ݬ��������b)Z�֬��v3������YU?_�?�qU.��y?��WX�ض��t{�p?ĽJB��м�Qkˤ~[h��f��ٺ�֝����tT���K����S޶2yѕȏ��}'R̐C4A�p��|.�B�Oh��Sv�f�����-΢\"�*�����}��_�{��M}97>��;\�э�*_�U����d�Wl�A�C\��29��Φ�k��r�WB���X���al��2����&Z@�vE�y���;���7��dM܊��c�In��^q���6��^ێig����yrS�:���4�KG@���{�E�A}˯G��Dy䌛h��n��m���vX��Y���Ns ��/�(�����z�'un�'����2x��{���L���m[|Y����5WqE���~U�i�kjp��Z��j�(���\����@�p�b���~r�:�%[�V��k69"��kH�E�z�^5��鼢UİG�"��&<鋜Fo>I��q�U�a��tt�i)�(�����+�~���f)l��$>���n�X����ΰL�����c��H-�Y��t�#���ظa��\��r`��&�p�Y\���-_h����
����e�x�O��6=u�8�~�8[��j��Q�x���>��að7xj\��X ��_0@��(>�$-?�n{WUw�,*(/�6��ι���	��s._L�g�9m�ȑ�zFO H8��?�};>�k��Lrn�k�	�bm�Ε�8�5��w��Y+��:d�{Z�@�p�]/�x�;ЊҬ�r�i�t������ȸ�� ���(����G�k�m�l��&����. q
A�%�p�A�TbKv ���Ed��Fh�eG���F}�U˺}��xP���5У�][�Y��{��A�y�ݖ��7 �f��uخ��v��nn��.n(��cq��G�vr!�������o�����:O�?�#ި@3�B�G���/��wp�9ѵ�
�u4��<Z.�����G�[��k�v���8%��p,�怆t�\	�+!���ā�)j��d8|m�"C���#'S�xR�u6�9N�د|u�V6��F���6��֑*��Ū0�(�mЀA7�0�@�\�[_5V�Y�K"2�XY�A7wж�	��_��J���B�����S'�'�0v&n:���pujAa��#���eZ��{��L+�/8�:�?����b��lѡ��½Z�#��z5j�˔i�����j3ؕZ*�@/J��lr!�}�O���I��J�O��O6�)	����F� ��a�fB�U�W`�wWN2��&���ь����F����ܑ��`�e.��̿��H�<B�m�`�{b��7�4����"Ũ�Ǎ+������
���q5����ڇ��є	�)o-�� �\Q�v�+�?'�Q�p���u�����K���W����u��.��W�[Pk�*����(=ٸ�"
�Q7p�m|���TH�~E]_�jyqA|Xj3��h�r�����W�ɞ��?t?�e~,��j�i�?���\�L0����w<<^��6t(�3h���)-�:�ئ�N�8r	��!��#dn�?^�}��^R��ܰgφ����h���  Y���AX�X?6*����o*���)K�>���H���<\���M���)G\k^�N�Q���w�o�#q��wB�
�l4�T�p ���U=����sUH�:Ֆ��?���S�ͭ��j�ɻQ�}����i�m��G�B?D����7z�2�h���{�62QNߌ�i c`�W�CYJ-^�Y�Cg9��8}[49����K�w<ꔕ)%|}��+��)!հ�?Gь�qU��(%��rۆ�)�R5ko��S�b G���k��+f��M��uY���s�23D�nR8�I�� �X��+��Iɑ�'�]�
���u�8��jة@�3l=��-k{�-�hg�&�ѵLLF��20~��
�4ծ�43і�����ɭ#z�Ӆ���!���7`�K�ɦ�ٝ�\���~�"u����V�,��*n�]��}��^��#�߯�M�w7Hϙ"����Na
c@� ]�#˷�����.ƚ��@�36��'xx������w��A�S�:x����o&L���Y=���	��03ʏD�3�*tE��)��?�REY��1�k�Oi�k,Ф����mȕ/8�E�U�~ˇ�j�����e��K{�2,|��k%e��)�</k����!^^͢�4nG:s;,V7�*��|�m{z��4�[qڊ]�*�5�BO|�	d�;ד��>�d�t��D���Sݱ���ܬ��O2��mLn�� ��Ct���M���b �r�D����~i�(K�S�.��Ж��:��`�w�[��p��������ah$�T���B��D'/�^��Ce`�C�)ֽ�Ch5,�;e-���tT�;Zqd�I�-��Fs��9�|m#�­w�`�6�1�������i-�$J�A h�jN������h�u�C+?;���$2�.���9�s� ���v㌘�Q`|��������8��ݪĸ�`D{��n�*^ͤS�7=�]�@1,�!��+7�|L�k"K�L
8�p�S6H3$ׂ�O�#�m��v���
�+pk}Ec*܏��ۀeQ���ȍn��F��CP��|sF���ao���fD�����\��%Q�*�q�]�Yj�`#m���xr�7�.:�>�	]��
�� 	d��M�Jbt�������Z�4y��pUJge ���QϹ ���Hj�>�z}��L�ȗ�~J�J(��%��"$�(�L�<�
� �J� �cF�ǃ_!�lR��O�m�N�Cc�/�y� HH���%�3�O��*��$L�O�>�H*�$����&����*�)�5"_�tq%�1PZ2��\3��K`����Ho>�܊$���$?~�k�y��i~\�9�ԯ�eƴ�U��QD_�/b��J.K���:��᳏y��-"��Z\�5®t[hvp��c"tN@!<��l����@�����T?W���̐)FIL(�:���M�m5>L=���@�ިU�VCK�y��	m��T�=��"��U���+�t��(T4�ū��V��A�㜻�	Aܱ�wM��/T: ��Xf��;����,�؇�B���Ah$K�=�V��d��l�	;�L�
RA�`7
d5���s�"B~��}
�L"q|��' �<�#��f-�ӎ������33݉~}A��ڈ� �F� ?�YQ���!�5�r�"��cmg�-m���Ȭ���+��u�=�f��<�ͅq[Sk�;8I�yv���ɯf����5�q IG���G�`�}�� �����yV�Ϳ�Χ��������01�&K�Q�����?�[��ۓWE#�t����j�k_đg�&�M��ӧU�Y���A��Q{n�!�"B��?V��y�$� �]6=�
>K�yנ��~PF�*�4���f|w������­ 5��s��C1]�� T%\��uW7�zP�FVcJ���!���;�\�_/3J��H��ߏ6�DNς�:�#ģ�Ɵ�Il3vbGP���QL7kn%��(�J����H,=�	ܹ/��9�:S�����hNP�`ӔS��-�+\Г�:-c�Z7��`_F 9��z���ƬN4ElV��AIl"i�G'��y!V#�ݥ6x��G�����%�~R�6�:n@t��Z��g���if�X�ј�i�qv`��y$<�!�*���ԛU�!�-Y�p��Oڹk'+M���8��0�����L
��	x�+�{f����h���.1ԣ��-+���=������G�� �ؾ�{A ^�/�e��"%U��R$��O��6�t(�� ���z�A�ղ �����`,����4l �"�olvr)V���C��Mۘ?k嫎��ɴ�2	K$ۇV�lϙP���[�p��W��k�|Te,��,�%������JbcF�3vۈY��t�tS,A��#ō�O�9��4c�0��i�*[t��RM��!�j]_!48h�lD���5�2aS�@<fn��f
���߇�0A8��>�� V�'�^��S��Q��k����m<G�F6�%�T4�i����W��BڶP��R�JpA����J*�OC��L�|Aj���k*�����2ϜȺ��Z��DN���	�ҹ�L�-�Y��T=�Y���͹�����?'5��O��[���zALV��G6��H�jG�o/������9�@ ��Ym�����(�
[��b&YH�3s@�]�N�*�an@��<����M3�p�vk��w���PĸK!CC��ڨDF��Y|�H�W����*��/��L�N&��y�i����+d�O�f��b����ñy2m�Y���"��5�(����&�{|����H�h7��I�Տ��M�s��H���<�8jȴL��'޾�ٽa�G�=㶺yv�E|�^�*�$5Z�
G\��eϪ�Z�|���[9k�U,�-0q"
�Yg�.&��|�,��%��S�b�ݼ��[��^�>Q��&RV���4���?a��s����!<���\��E�sO��[J��N�;����,3������{��l�u�t����#f��C��Ci4�ݰ�(|:�b��ԩM�eS�^��I�ֲ[��X|4�Ї�Eg7�ݴE�y�骋|S�#���]~��\���>��� Y��F��iI:f��i-�aE&�#�J��3���y���}ݙ|����
�� ���tb��YZHM�"��N�[Ԧ��@P�b��|���\�@�஼�n���xle�=	����S;�[)��y��?#���˪�M<^����';�`Ơ��W��o��H�1�f�ư{r����Ʈ�J���!����+��²��|k����eh����ol.e�h��bCб;�kFgh���#�,8��8�^p}@*b�ל����7�0�]y��.�%�
���2���Yd00��*��/�ò�f z��b;�F��Yߧ"�T;l5
3O�h��d��V?�?����>�"�P.�ަ�������O��CK�G�3kf/g�[�L}�/�׾]�3�Q�eDl<9I&�q�"�g��������3�82ր������#q����v���}̔x�0J�k����pm��x�Gv/��9��b���K�|�(g�M2�4�Q�.� �?���)��Ɣ)��5Ŕb"�5r"&�v��I�� ���J���/�7�%�!`3O����:�=�MBq8P#��Q��{n.gԸ��f���mǇ�w=�r����w�Ј���(���Mhu�l�u:�=LM�u!�i,�tS��N��&��z$�+OG�&�X-փ(� :�?�����'W*y@��E�jk�n���R�-�MK@2�4g.]�,��J"_�G����>Vɳ��\��.��S'�i�����Xg�D�v:�7�޾�㽶�*����/�n�b�Q�Q�C��`Xx)������������tQ�\@	>J�dh��J ���<h,�ԛ��O�J�쏶M���՚�먳�d��Q��996 �Z~�Rl����#�ʓ����޺29w���,�φ�����3?V���}f l��.܆!����6ҀSv���1����[.bC��q���e��������zծ�?u]�d��}�7�{w*c��9ꗁ�[������d"vW�|�G����K�������jB	c`�!0r�o�6wW�y�j�7���/>1R0�L)��<B��K����V9��N"P�Az�R����� Om���3ya��:[*����_��_�����=g?�<8��a����#-&�_�b6�)�r��ܣ�3�\�P�d@䢽=S�\��Kk y"�����ޡ�����9�����ۀ�z�����"e�Q=r[l��K/����&!y�f�O֍���1�G˥ˣ�-�M������z1s�^}hp�����dTw���x�-XTC���n��)��T)��*�� [o`�t�K������ɵ,���4W�5w]tc����g{ l=�r��z��J�xF�;@�6H�Tk��,����V�:p�z����2�& �|�i�aZ��'F��4�p[�A�G8jJ����ټ�Կ�}<�d_���U������S��3²͵V�miS�kL�\��W2/~U/ŋ|H��& �R����*��0���DvV�MG�L��-��,*��`~�Y�L�ڎ���3_�jג�!a�
D�'������=.��@,&xd���I]�l �[��t�b/3k����L	nb�E~�Ӏ�� a���٣��I��3<�d�S�߰���m���&WG��e��_�W����l�&|��Ϩ�,�C����>\(�phR}&�p
w�#���U+��7Ҕ%x~��:��M��9e�����ч\z�]�%��0����9����/��bN��i5�L#x��wH,/�+0�]�v��˰~���ug����G�z�M71o1�S��xqi?�j�
�Qz��&\�>jk�D����[��O�c�ja�=�ȉ�<~`=�x�a�Q�p����P�u"kyt=Z�w�,�]5E���	S�ȃ4JɁ��W�P(&j�V�D�OT�}�� _�S�X�F+rCAC%h_8֖�(��W�O�@z��)k$9�\=0���J�����f����2~m�f�*��i@]����o����"B�$Vݧ��B�Ld�P�FhQ뿎G �_��\*�-��S�Z8	�9)�����{�5|HC!M� I:�ݳ�Y�����%���=��3��k����O�_����\̈��1�� �ʥD>��;-�ҥ��߲;���:Y$iqqJq��1�3�w��.J{�sb|(t�Ln*I��wu{I�~��L�[)65�:��F�9q��5�6������O����D���z�t8���б�/yI5L�:Z�_=W���А�RҴ�7i�Dn��K�x��S�,�e�Y�E��ӵe|m��� U�)E�!Gy(��Xx6��c�_������M5Zm�H�#��(����
HqNk����g���2�8 ��V]��9R�q�O��T}\EO-��b�뾮���O����w���|#�{E�s��r�鐘$����d\g=�O�*�e���g��X�?����Ė>ck�O߅w	X���� %!�k½z�q9���(-E����ica��H{,.�|���p/�t$'G.�*��!�qR����/�A3�r�v�lہ�����$ڗE,#Āf9�-����xj�O�&�L���n�����(!��Ѫ{E
��dq�B���8OX,uY��W�m������*&'���bSIb�pc=u{�%y�B�#���^-�)��Ȇ���m߇������F��,aL9��`94��&��i^�E۴�H��������{L�;@j<Yhx��q�DӫL]kd�ͬ䋓?����7�atX����QT�������0��~�	8�9c�ב��u���c�=��X�^�B
P?@��&X��B����t�H5Ɂ��^E���:p�t��99�|a;3�N���+�r_�*���˱U�#��k1?�8n��c,��L��bBG0�:߾�'#st�� �/��oz�RAK�P�Ǐ�e.���fձ2�bX�-�:v�ힼ�"�X9-mӽ���βz�ì��	G�����,���&���8��^����b�F%�:~BAO>��D]��$)Dv��
_�&�q�Ww9�C�Zuh���XB��k@�A2*R�;7�B�DL�m�e�?<�؉;�cPƆ��MQ���Wx}Ȝ�=0��A �=������1V��Ϊ�K�WP$�RR�����W`WqF�2��c��%ǵ�-��-Xs�kǠ��F\��9�e^�����翖��]���<n���������<�6+�<�"��?nT0/L@IM�]c��1�ES�^�� .O`��c)r��1�0�'��P��]��](f@�����3�(���&����BbJ19�Tc1u�M�Z�� >�f>�ԭЃt����,;���\��s�a���%��0O"�݊���(,
��7�rdc����2OQ�K	rp��"���n��l�؞��c�q�e�k�~~�A:Ml�=[v �He�ECx��J���Y�Pޓ%�w#�
R�wW�A��%��E�)��I�sD�]r��q'�E����S�cE��y�{��ܾ�q�C����#xl���-
�җ��*%�����n�֫#�Ǡ0'�w]��
���8U��-:U��� ��RPǟ8�H���哌�$V�8vN0�L�߮��tfo��z&�
�ҋ2�5��d��Ɛ7ٳ����xd�w�R)-��F� aIq������u~�&ER{i�p�τSp�j-�Ϭ�p6�}�=bY��ٹpp��F�U��3���������v^����vT��S�<�?�=���1�7vA��^�@���.���ڞ}�iG$�Vhؕo��v��$�w�qÐ�g����a�ؼg�N��/�)�׉~��Y�:�q�L���b�a4y��O�(����2�"�u�l��Z�.,����b0�x�8����*�ԫL�kN���F�c�\��/��q��|���,�C���,u�idis+�����̔�7XT�oU��({r\Zy!W����o�*�~h�D��Uhq�- �XW$�k�2]L�2�.1E0&���g��Qw2��낷�gg�Q��7�����6��)x!�X=�]��2r@�OF�kɄژԽU�-{�����1ˌp�����u%��!�}=e�B�%�`|��_��+T��#	�7ȓ39u�;�yDc�E���2���L`�V�e ���Ѩ��q�L���V�S�6ug(�G$h���q~�K,�_�F�V,�]Ỏ�Bb��^���>��;�T`W��TCqEn9`tHm��̔e`�ه�I봔�㩚���A��w�췓
w�Dsm��R�U`~=2U�G�6���[5�u5�s"]�
v��;���xv�*���w:d��),V�m��4D����ހ9�@H�6f<��Ueq�������u1EϱH]'�ȍ_d��6��:E
M��/��6�3ln�=��լ�n����D��5��|�Q�>jO�MAx��G�F�����0-��� �����I��U-WU�$�J������|�����a607��b�э�pF
��@�v!��( d�6m,K�t4Z��l�zFl\����5��+x+蒬�F�7� ~É����kr�MjRbR�1�rW��d�_x�y������B��_͒^�Y�#SyA���o�JK����Bͧ�uL.�|/�Ei,������m�Я�[p-�9����	�B�_Bεl��O��m��d����F4k�g����ϋ0>_����}zo����*:�Բ���u�>�s7[��B�ʋ���pM�1vV�H����� �Yzz`	�r�X�?+�^�~���F�/�7��Af��N%��*H��͈���k�Ȇ@k�M*�'����{�����C�,C����
�OgH5�#ݹB���HN���0S˚O������<g#�+�Kox	�ޡfo���MVuƜvK���p@R���;4u��Wjy�BO�w�`Y��Ul�Y��I2d�A#��s�ק�Q]Am��7w��/-�_�H1�L��wi}�Ï�y�kVq�I7��n��c��4��_yuu���(\x�n�A`����3i�wՍE�5�#~�3��q,�ۄ�JS�]���"�A]p����YmR��(�堁/UD����ت�!�ʮUW̼N�3���)r� �q)���x��=��������H�nk�����G`�n�
�>�:����`���~�%�+�'p.[����Eez���2P@�E�,��3ࠈ����K��nZ�u�Ps��+��W@g�cL�>8�8�?0$e`=�d��O5+^���v�	F0���T~O@t�C��2�Bܿ�;�C�r-�J*����0#�$�#�9�,� 
.�l�$I���Li��z�tg��芤i`ܒ�P�W�&�lrwve�b;�d�r�$��m��-��&�����Ǒ;��T"
޹X�ys��K�������a#���O�[�O�Y��rsX�j�EK� _��G��w/�-�Z� Ƭ1	�Q�M��ARιI9�mԙ���;��m�ښ��2�������=� 	8wz<y��zƳ����rt>4��ho�Des�0CE����Vc�n�	f�E�p�ޅv+�+��̖K8;f�6���m,Ћ7@�im������f�T]�'^��P���bg�˵�*�,�8��A痄ߠ��q%�+��3H8Nr�S��[	z�{;ǿ�a��ہq�g��L����W��n��s�I.���46ru�Xл6CK̴ih�E�!T
����p���V<��8�e��_��Ø�1UdN��ÜL�c
{5LU�O�����?�)i6�۟�FM�����?��B�b��D�W���yZ���)��-VtO���bu	�#�f�:�x�H���A�-�\t?)k܍�E\��4�@�Ex�����=�L�3��6/�1�Bw5}����U�]�f,���k�����qL�>�q'�(�������TS��3�9�ڱ��_iV�a>�
7N���bJN�\�|�b]�����~y�H���IA�|�:�s9]zb)�W�_��taXao�`�����`Ա콻+��Kݓ;$�J��.�Z�5WZ��=�.>\�'r��vx������a�Ճ��#�A$1�X�Qz�((���Z��s0�$!��)�Y���[�	]��k�4���"+lx�B"f�RSX�o��v��&D�_�.����[��V9�L��ԡM��*��q�[�%����8�ߛ!E�G�|� <�U��$8q¸�x�!�18��~��X��2��ږ���]1ZL�
9�X�f<�����v���w�b�C_P|��n�Α���aSl�HZ���T�vm���ل�ޟ�8S�(�ˀ�dQ`͙#��L�"k�� .�.�/g	;�{t���eT����F����~�m_;b䜧����ϙ�8��p�"�P'�Y�h�`�} $2}W�bE���I94�)������͞����G|d�?xbN��0�i�澣;Tw}�<F>�mwx�7��|�&2�=}�0�2[�9�._�f��`9�W|F>@u6�̎��c"�#�>A�1�G" ;if�*N��f-���U�x�v���[�����4�Y"�1�΀SgBQ	r'l����F�!�c�		C�#oy�Lͤi���4KcBٿ��QZ5 �j�q��=����n����jC0�Ug��t�_b��ǈ�Q���^H6aUH����X��3P��&V9�ȟ���z�z�m��]���ɗU���t����YȊf�=���� h@1��o����b +�s)X�B$�|\h!�fv�lvs�'E��	����ND3,)�xd"�VY�hy����b��'��%�I�o;�y�spOlu;�)�)�[:JK&�ڿ�܋�O [�0?�+��/j&�x9 ĉ��כC�Ol-�~(<2�gG��O��Nʆ-W�}W�4^���[�� ������acL/-r��a��*���1��"E%HWb����,�R����K^�/���B�`mɸO�T�y!Z�#�&�ɤ�dz��b��/:�2j�4�A���=O�&�,�����W��9*���B��ֶ)΄<�b�ˁ
J����8�^���F@���`�	)�B������
c��MY_Vߠ���������V);(��{O��T(.kMOO�n�.��a6s|M�=Z�2�N=!�O�SIbR-D4V�������h�\P�ؽId0-Z�Ne�C�	I����w� ��X������L
ja�0����y��E=�M�Cт�H�#�{`8�"����Ff�K_�W,j��w1ڟ� ;���$��Vw���]�G�U��FQ�oS {>K�S�+��j�z��\1�#[J�3E���b�J��ܪe�K������)��q�a��ǶILw�׆ <F�,2���!�_@_��a���e(o�+Ed���(W�dz$"r��[&��F;-i��d�����	��X�&�h������%���(y4�
�8w������m2Xd�|���(x�D��۬֓:�1H_��u)�Ǜ�\��uf��D�����S��.[�7���C<B�^�^��g��K�;o���* XTv��<9:���%��1��hL�5�����ltI�)UDC���5�]��.�B��}�鮊	��1N&��G���PT�o��}4#�+j�HV=�ǻ��!|�E��.ӵ�|<@�A�D-�5$�jN�	�&7_�ßD��рS�U��`���C���!2Q�>�[�ӥ_��^BW�_���ғ�AH��a(��LW9-���0�^d@v	^��ݙ��>���X�Fj�N|��N�&��^��噟}7�������j�0��8�֔,d�͢T��(�nd�����q���!�P`b�t��~sG���
����w�oA��`�
��U���i��ZgP�8.�����JLP�RɐrIC*W�Hc�+�;^�� %�f_)i!b�\K0�����l��*����8���������ض�˺A,����Y��)�^�>�H*~��	����H�D�����D���7�8۴�q\��Y`���ζ���w�Drf�˱���Q]F���먻��K~����?���@�u�yr�^FL����4N���r��u�<��\��v����Gu�28$�?6��'�$�@��r�x�8�&9�jPx�����J%�b"[�+,�d��ˡ6�)j>�5����E~�C�ڋ��	|N�%ԉ��{�_�r�2��j�i�g܋7�a|([#�k� ���Q��,p$��ۦ��W ���<���	����w���l�3��ԭw�#_��\1:�bmھ��9��B�	��@�8�]�u���S��#R}�$;���gI���� G˝fןz�p0��+���C�?@������Dy���pU9�Q}�=B����j-�ŎhVP��5���}�(Q�G��c�;u�,۵�B\\�B�k�1Þ�x�6�>u3>ɟa��|��
g���%ݩmY�0�����,���D)�X�w���O�$��f@:��Gø^)��H��,n��m���,I���E,��u�6�����׻q�7)V�{6튱(�_][��2��EC�)�D����sB��v�:#�_|B�����2�o.S��zT���/�(���d;$o�GᏩ���vmnI�r�m60�_ i�!q��� �E{�?R	��i�[�]^t �ґS�}وmu�����Q�7����ǂ�k5=[���������h��D�Y�]��~\�YO�M��~��J�<�k��}bq��I~�����Y\Q��\"Å�m�p$�q���(X�>�Jn�X��IP��lC��Ò��u�,��hd�aws>�m���|l�_�~_����͗��ڔ�s�`�U�!`!l�̠��!K㦱��v'��}Ӈ獑<����1�L�m,�W@r�	 uhMԼ�W�I�ݹ��j�>� �y��s6i��{p	��rPK{fs׿x�1{�nP��ƤG��S����,J�R��RK������i�0�*9ՇR ����I��$��p�z/�
�a��Z46��Yտ��Da&�ژ�s�N��ME'V�z�̠	���EF_b2�%&�B絟�|A���JE��M2K4ן[� �EE��o�#h���f�tP}��Q5�
�3,�\�;�f�������r���.�Lv���ۆ�a�|��Q��(��G�a���P�뻧��HI�|c�Y�:�gC����lYk�vu�$��/�zh���`~��O�Șm��;�k�Vo�QG0W�XK��x�hy��jmD�+%#II��MDp��p�;�(T�<���0�	#�Fq�E�$wML���=X$O�G���e*�iK���6�3�JG�=�6͢��+�	{}xp1�lDe`���q�B�E���1���2A@n$���\�Ө�t��N�\�Y[`��#On���2t��d2�_%b� ꀋL+��ӧ A���h�}��y�� �$��H�oj����J6���cBl'�(0�Y����/֑�G��pg&�]	�Ҫe�{�ԕ)�QƳ� ��a�d��]" �]� Օ�I�3���W�b"/��ʣn�~�$�Y�BG�H҇�����B����	��c��C6��f��;Iq�Z�٩q��_=�j`S'7�e���,x*f�Y<�f�]*�?�b�����徘nt��=�ɸ��$0�Y�K��R�]D��B\�o����Zj�u��E4�,��k����v �A}(�q�:c�å�eɋ��������D�\���� f-���J��-4�DT����S�=C�s-,2V��(
��w�^7�v�k��:�%�J��(y���{�jH6,�6�:�T7��{�ԲD��p���W� 5���,Ith;�B���+�uQ0��R�:�H�-4W��߹����E&�R�����N6�\�������(H�f����EZG�L!����_#X��L0��C
gژ�Y�W�r",���1�"�Ć�c����}[�7%:| �������Hz_]/�嗨\	¿!l�U<7u�.~��)~{�=Ĉ߻��ޖ�Y[���B�T`-�$ĵ��+�V� ,4��[NUT]=o{�R
→�*�u���J����vH���H\O�)m8A )��u�fUҳY�1+ �8�Ŝe�sPv��v������~�&0��C�X�ׇGG�"���"�Bω�Q~���n�ƉI�a�5_��w;k��
e�l�'J��|���>ya�ф���DR�h�R� ��>tm{����?����Sf���λp-��_j+C��S���S_�	P�_��n�Q[p���De��1�u����
���/>b�Hj�2}��Ͼ�L�+������7�]�*%�M����������h��B��G�F�����I����or`<�,�;��'z�˄�|,�4@_J<ŋk�%=���k�o�A��]0������%�P�͢�w7X�Ci�ɼ��p2[�46<�sgզ4�@6]�y�Mk�r4<В�M�3M'�4�ý I���
;�м+3�C�ߑ�)M�L���v����'x%��g��[�$����Vj�&�<%A"�Oq7�CzA�3�z]�zɹ�*�y��7�P��)Xtc�h�����d���}���m�a����EZD��D�|��8�m-3��6�c���-I&|��	i
r��AM�	�w���f����8��`
D��)����j.��8)����X�U�G��4e��·.S\�� L��(������T_��x#Mϳ�v�]������_�zx��4L9L���̴B2�w%c�߮�c+a�}c�U���;�C�`"��p�~O�V���S��F����O����c�y1���ߓ뗩���9���e!��>��y�: ��O�����3�����D�R �=<�]�IT,�Y��J8V$��o%q}�[H��*�Y
yv�/��Gp�#�%�7x4?��|��������W���6��J2<�/e�Y�-`��cjXH��b�&�e~�K�H=o�.8IHL����)��̾b�i� ��������B�	�1.��ܯ�t�`0�%��~K1A�/[]$�R�����>c�L���W�D�=*#�?^�sGF}e��:��WY�᢮~�vC�eT���ꪄn�$G[��{�oA`��Z�e�Z�ͫ��p�fD^�ڮ�� ��7� Ye���(Y#�AAr�
�
�m\��8wn�R�š��ݱ�-����MI}�=��G,N%�D=O�ůk��c_�g
�u�@*�|n�� 4G��e����� ����QJP��RFn}a�% �QQ5,Tã|�����A�L��?�J.��Gx(<�BUx*\Tӫ$8ca��f�k�D�z@9��^ӹ)�%����Ɵ!�UTG���ٰ�|���a�����w��g��
��inA{6�bc�fx� �V�F����7�+�F��zA[�y�i����S�RQ_.�92�ȧ�H	6����#���}��<��m�.�[�j���ٰ�T�xu��o���K�jDk	ي�������Dse�`�t�r�p��L���ql�>IR2����k6X����DVceO�����}�?i2U>���2�'�T�~i�nHĈ��,*g291��A�_XX�2�;ɛ�����~&4b {4w�������R÷�����0B�6f|7�U�=��~^���_�"h^>�Ih������N�B^7�@�������FǢ�?%���j�P3�5E�1�O�o��
�瑦:J����}���zV���Z�WT+Չ����#��ş��j�7s�;V@�4,���ٟ�����)�
ZL<~�?O��(L�ߒN�c$�M�{�KWne-��2�z��ė�������ݮfi"��l!)�@��r:�&��z�d�x�tL�p��/�T,�f8(!��לC�Ecv�֏"<�w{��K�����x��B��1�:���;�_�t~�"@���o���+N�\~! Y����i��b\���QL�)#�cБ��Wߙ`|��y��	Q ��^���^r�P$i�U�Y��B�v��[�P�g7�IE��) �O�iʊ)y#7$��U�y���o�z��5Q��?��}�R�B���(�F�p�����f̹Zew�!�D�)���-�n}t��lg��j:6�7�<}���v`u�'0�\�k�o��"������,���+����Bg�gp�@�E$�&SZ�NY
 ����Y����v%���_<C��H��i�?��w��R����sz�.�
@f�;�1�?�R�S�Ђ6�����Ͽ.x��?U���I�Q��'Ϩh��.�����?�Ho�Q�3�xF�b(� �%eTV#a{6��R�P;����_�C�¼�Ǝ�Q �������������+��p���̢��`E3.��;��*�4�_
ߘhN���Q )��<�]�����́ I�k'$��E5t;�	�V�1�A��T�liV\gƠY�{�F;3��A����n.Ŵ�Y�ZF<+p���i��сk�H�gy��i �x����Őz�Bǥc����?2�M C�(�� "Մ[�},�`��Ν��X}��=�J�w�7�w�KF�sbKx�K��Lr$�8n���=�AF�����Qy��!�WK�o�|Hä��+�+)��?��%�J5��-��$	I{�MbA�D�ʰYE��-��ϨH������վ��c#��`��SI�S�p�Λ����h�z����>$����|��@B���u+�6�[�k:ρ(�������N`!�Gv�^����'f��l�iR,��p��cl��(�
�O%���m�&��=�Ż������G��L�S|�������!���l�M���G-o?�E��eo�V<��X��,��������,����O�"�#���c�[.�M�H�ƩH��x������'�s'lO��~~�g���}F�'tu����Ah��F ��~�~�`�<�/H��,�k�H��ߏ[T���c�EM9��@I��-ä$��~U�K�	� ����H�)�h��N�a�+*��N����y�(�Ul�E�%E���9mSך8��m�����sTq"�����6 o8}:���j�-Stz��sR�ؗKnL'	�=�na\�{-���S�̢⪻[�dQg���t�;�&ҝ���[��/OHׯ��1z�;��d���8$��I��؝+ E�v��@M'W>��?\��\����d�z/{���?Z���:���d���0�����^!5|�r�+�_8Á@���?�i(U�:�ڏ�;����Jy���p������i'h�:��Q�A���V8�tU$��ֻ��L��,A��"D�E���"���z�&:dp�IJ&��i�iC����'��j5��R���R(���K� �e�A�����1�W�pha����>�)SEq�e��"�Zq�u�$C��;%e��#	�P��]���[��`nS���:ؗ߰����e%qV��e�R3 K2(��:0�I�KC�����1\��W;u"�)��c�}���xb.Ai�L(Xa�����|+$R9��	?F��~�	�T^XX�h�L��΋\w�n(W&"��N�n� ���5�W����pO�h�4�����5��0���1�[=Q��5#3�e�}��~���'�I��͙T��FByFcD�Lz6��,侩e�ЮPV}x���	=fiN�8��g�y��S��H���f���Vت[{ĸ��&X>O��>R+�	���
�T2����P��:4#���"g�������/26�����5�Z��i_b��,�L�.U��_,q���ksOg��g��m���"d܍�ӣ�^WaW0���J��s������_LJ�2�6�n\W�}jH��wn����f�e��c��������4�#�k����@�u�p�5��Z8�T-�W�s}��W�h}���ntH�9Gu�IW�p��pP��O�:� �X)�_��F��@���B���Zt��6I���n3$��A�[JI��6^'�]s��C�w��SS=9�gf��5�S��������� ���IR��wOB6t+�<���a�<���}��B(�����ç7�[��҅�����&*vwd����P����ic4fd����,	dW������}�����;�m�Z��ڱA���ڡ�ft��2(�h�;�d<4�2|@���r�8N��z����h5��~`���[�6k�<�v뺘����ٴ���Uy��;һ����xq���a�ku�TP
��*�������V�};�r\J��[%'@�:�+d��C��Wwz:`��?W����%����E�ӿ�}ك�2ԪLFe��r	P^	ʅHm�J��w��K��B��đ8��k8o':JK�����W�dS��x�LT��c��D�>O陜H5�<���J����2���驰����V�߶�jI?��C�x#�"�e5����סW �J^\ ��A��x_�����S��h4"���⎓�l4�A�C�d�F<5^�+41B�&�w^m[3Q�{2��8o7o��8�d$�7�Y�w>"+ѓ������/
y�����ǳ��:�1�� l���ǅp�����St,=v�8��@!-x-T��UC����ïKX�}�sb@n�S����-GECWs{!�N��7<Ժə.��D�n���5�mĜc���HJ#�U����2�9�|]F��>F���|eo�oL�]��d&�Q��ûKO��0S
��S�����:�d��X�Lҗ5X�K>���	'a����PM8�x�}Y6b^{���[�W��d�Dْݘ�V P�.�v}��5�O���X�V*#�la
�/Rx���ށ#�3�l�k�����+?���|J���7֏z}3����U��Ra|��gl�>�M����\�f�^o-�����,��RVh/�����W���I`��=7� f���7�^!��/����qf�s����#�e���2������b�%s���-�y���q'_tF�m�L[$�g�$��3������`��j1ڈ��p��m����!q�ꓤebc�%��7�':�� 9�W ��$�S�0.Y]d7���7��,J0��-U�0���(���pkiiǬabFj�^BO]_HbpS@�Į��SA�������J^�~�}I\�O)$!��T��̳�ߠ�l��o*KGfe��x�;�n�C�����/��{�:��.I���nz�����-:]A�	_�#1�7*����D�pr3vۑ����n�g��A3�fm�a�����+>�Xg�b���䗭A�D���������1;���=J�ci���ߵ���h�ː4���<����i���- 'Ƽ�Ky�%/p~�71��B�B�����t�a!Ā�G˟d����|��GT:7�1K�$��Ң�8Y��Xl�##�*��w����~�0b��5�j�����պ3�H �b�0K%��HJƅŜ����G��T�y�%_b���մ�>�yZ�.�N�Q�;{=<f�5���538%����|�0C��m&�c�|�}���K�l'�̃��/M��n�ޱ504�N�\��p`ة���G}��:��9Y��Hr����X��.p�/c09V�;���Frw��� M1��*���&��:�9I�}��z֖����*���]��fa�|ZLIƪ��r�q��+ʐ:��Ô��W�ƍH���ha?�r�^�X��U�#��{x#�62p������>$�.^� 2��8��1~��k!NST��lm��+�A:	!���8^LB����^�r�ا�?�nr�v�`|ѷ�;�@,����1C��b�@��H�/S���x�;����4;ܟ|�!���q�9�?��12��됩S���/<V"�h�����<J_�
��>^��d�m���>�zX�=6u����g� ┯�'1���HU��~"�=�a�+䈔�����`;N��r0M`���ռv'y63��``����;(����!
Yj	�]Vn�����!��j����9\��.t�k+v!��9-���T�3 ��Qr���u�"��V���{�wM��܅x0v
��0�A���W1����D��c�%ͨ�����
h�-�rV=k*�$h�8�I)��;+�\V2x*�bN������VD�6���%��e�AN�VY�8�g�l�|�a�-�RW����YP�>L�M��>k�A��*ȗn2�kK�N0a㟐8��{�]A���S�~��p�N7����9%���]$�2�lU�$V��FJ�JA��f�vc��rkR��8�t�(�.�ė(t�Y@x��֌�h/��8a[��E{�ɐ�4�%w��A��K�n��ߚ*?���+c���S�B~���dT� ��|~�L��M��Ω�~MtE��#}�Q�G�ɶ�����ѳ�"��&�;˸J�Q���bu*��UI%�b5ڈ�L�8�I��\]��
�A}���IQ~W��=�9��>�_=2VA���:��7� ��N[E]�G%}іz�ؒ8xXi�<���;�(>N�$�:B����V_�Ѓz��Tv���?yb	xeW�8�^%K��������P�7���И���3�ʨr։����Q���x�=��e���ˈ��/�BjQkӢ��E�J���_�Nb�V����~@��ٺ� /�#J���K
u�|�^�t�\�IK�V�g�Jh[�Dg��YzK^�9�5��}��=̩x=M]�ͬ4EG\a�hb��[u��J���s�$��5a�d��䯛�H�����ד$ ��]���x����������튥��a�	͒�]�1��XaR1MR�E�S4ˏQ����S|'	�р&Qǀ����Ք���녃a��^�,g��� Ucu�ͽ�{ɽ�����5��.��<�.잗�s�7��~�m=>@;�x�;M$E\:����zao��J��_(��ԣ=/����@wA�>�`E�v𣏕C����8�� �
0��mg�*�hUZ�̵f;�_O��s����\�\��?@��%���Z��� ����%�З=�\��'�s'7A9h)��o��']5�1�D�^-���١��~�r�7@;�}pV�e'���\'_N�sIK����1��.��p"RY}�Ƹ�&:�����EN��zj���#���3�yK/�Bq�����Rj�Dm�I]�L�#x���M%'�˽�L&�VK��	8�V��J��Am[U.��i�eR��Չ������jG��#��_���D��y��G`}���"�~]�?���� ���J�?~^b�nr�jh�Y��j��cq��܌t�trFM$�(��dW�ڨ2'���O5�����o�N[)T�8*�#juoB����IbxK{-��)!,6h����wL\yە�!��=6�4�F�u�h�,��{m�ɦv�75zI�z��������GS*�u�­���hx�ୂI��D��p�?x�S7xu�/?��{�yL��)p��o�Q� N^v$̀�y��M�q��wD��t�Q5�E���J�x:J��/o�c.ЧE)0��#�N�9�<��b�Jc�ÒB����P,����i��Ϯ�Jl"��'�������vՑ��=��T�Y�Hs�$����� ��5΀�7��:hi1�}-h�w^�4>ɳ��7q�\ӟl�y�%�ϟ��kX7�L��@s���$� �|&vi���؎N!}� ����;��d�t;���G�CF箧������b��[��ib&�X��n�5I�ј��& ��]�>n�)����B%ww�-�ҵ�*7� �����t����^b�hF�P��"Ypg�({�=%���V{�)���P�W�F�8�����@�M��4o����Mv��\ɰ��L�����rrP5���z
�WQ�؋^3DpDnN�6wܾ�9�7�@L��;�4�t6���[�z��+;=��I����)�97sY��G��p���vB��W�����r��w{�-��)c�j�j&	Y��G��
d�`�b`6��f��ۆb$Fę��Od�?G�u[~�e΄�z|�sЮ8�if��H�&|�[3����}w� ��[�t�J��Dv��oSQAK�/�=���66u�nJzq%R���W.�a��wq9�(�����7�)�b��'9�����%�턈~��aƤ9��'�3��_ݶ�0�^:/:�����f�����s �2��$0Mj�x	H�ѝ�ļ�	~��-���&�I���F$D�S��Z< D����2��m�T��C�t��Ʉ�Ʀ�3�6�+U�~L�������"���p��%u(���ڏ���!�
����W�U0<<��Λ��������?@����(+i�zO&	�g�B�sl�:�Y��7�f�������8��jTo7Hǚ��DS�I*�HA�̌,,(�ͳX��EE�(���/T���D�wkCC��+}��p1h���JP��\0��"��3:-��p�Ŧ���$Z*/��
���GN�ڸ��݅#�Y�`��S�����w�
و�\u~B��h�L��|����;�1t	�9Eݘ�)Q�-M�4��jݱ����Ԃ���`hspw0]�։����°[�T4���t�%F�BD��eǬ~��G�yǎAU �<>T���L���$(�yk�al�������H߶�	�b�\s��8��Bi�l�(�O�i���	p��g�-5�Rb�SFtk����;fr	���5ڴ̸Z|H������n*��VQ��Jy�x���P�~��1D�"���(���ruv}ޣ��%P^�����ff�>�g��z_��o��e��#=qq�`Y���3B���G:�ܴ�-�������iϣ__ͣX���_P�$���K�
ؓ���~�b_��b���!vj7'���V�;?��v `2/��3#ڽr���c6�ڔ� ��x��r�.���cRPٵ��s�����B>�h?�:��'r�S�}�#<��ʕʯ�P��!M�c�D�Tm��m�j�{��.xLqB������a�P���.ro[9��ƪ�N4���f�v`��ֿU�=յx-䊌7��+�(�����%Ux�G�(Y��#�v�E����U%�{Į�]zw�h���vIjJt�~��j��+�����.��N"f�:օ�7�'�[��]h&��sSr�p�5*�| 0�7ڕ�nX��{<�Nx�[�|�6�K�^B��3�~/N�+�u��e�k<Y4�+C{~�]�[Y]QI�#�;�N��&8���}'K%po�nڇ�C:�����f|H<?G��E���	ۦNe݁h���u\�ݚZ�#=�(M���9�^ ��0�@b�e�OuQ}6�-�l7�ƌ�@�	Ax�
#�(hT\�9��,1��ǟ�\�N�$�/�[�[I�B �+8P.�q��y�v��ʨ#���li�ȵ��b$���	���Y�`ѵU��
c+�V��)��H@��^�ݏ�6�{c��	|�(*�\6�����w=9���t�셄��>�|Nxd��A�.H&<ɉל�^�Hm�����=�,����tzs�g�6M��1��&�1C[��O���|I��i�Ix8$�'�p��ǘ�mJ,5�P>A����l9�h�`޹�@c�k>��*�d
�I�G���=N��B�V\h�0�M��\��3��a���%�j��°*��,C0�uͣ�1�m�;_O�幢.���>V\��ZPk��K�����(-�V�'��[@  *z�G?�m�Vs��+�Pt~M'���\�����3Qg���=v��11-'�4:	����O^�]���ĺ�a3�t�6����R�����:u�:� w��5s�g���ͫ�O����y��O���nW©�L��O�C�6�q@��x���j��W6)4=/M;�!�N%�L����tmB/�Ζb�<L������'�{.��{f�>$�<k,�����k۰�I;+�Vqt�u}Ҕ���ѱ]L�?�@ OUr~eU���"��Z?��i	|a���_X�6਒��u�KnW�$X�F��&�a$!��)a̯�6^��l�5�Bk�y�"�����ƑM>����,G��zVxz�m�I�(怙��]{�O�r���;D���;�7}�z�}`��)�Iwo���ם"���`�\�о�%��/�H�^�B.���a��9'�� G]2��8`��1�m� 5��-!���a��jJ�W��nEK�o��2�3���hA �n�!]Z��c����+:�Ԗ�z����hzGm&P��Y_W�&�� I����W���E��8]I;��T�ƌ�)R�� �`�^*��fLH[l�Jw�|����x�<0_�K�A��b��[ƙ3�HvK��D��͡#W���U�&H���M�}ru��P�]�#��/�������M�[��~�Ybg\q�D�k�n����)�"�5�A1٧�?\0,�h=]�;�����{�^ӟ����p)A����r!�VB��,�$F� ꆉ�5�W��t@C��bNJ}ζne,M�=Nm���K�C@d����p�p�6T�Yŗ՘��੶����A)����=��?�~(-OF�MCJ�� �	�#�*�-�e���I�`r49j�j":a5��Kˑ�\�MGmb�n�fl�O�̹��CG[�ٰ/}�?'�	�qŠ�r�N�x^��N�@EM� �T�a��)�Q҆���+�~	z�-��S�-�&<34�1݋?<&���F�\Z@��٠���ˑ�m#�GE�XGs1{����Y�T_0-���ǯ���$�?�c�S�nz��3�����%�(\�����R�{���f�ʮʦ�D[��P�hϢ�a�аߡ���LO)vMk�J��>V�K�66����Jj\E�m %�>��r񂖷D�G�նX{P<\B9Y�_�#�9dM����x���1�'
�@=C˗[��K��"~b�8\iJ?}�f>g$O&�_}+��B")��̉�(��-��c�i̹�`X�߱�/?v8�P�KR :�P�e���S�����h%q�vu�',����Y������^ �]e�R�q 1�>�_�6���V���Ȥ7-n#+�>�w�*�z��1C�F��U'���Z1�a���#N����к�H��S��_��䞸��� ��.���k��|��U��q(k@$�E�q%1/��Ss��4�Լw≬�,�w
��桅<�J~B^ǏR*E�5�i��9���G�����`5��������zU� e���
�²_�1�l������R�L4+,ʹ�M�^HKow�{�|�4�g��o[���8�c����nI�A��r؝��(���<\2U}W�nF�7�4�6ˬ8�-��.��C��1w&=���Ǟ���U�� �l	�ʈ/'���^��M��!�Og�4&�(��ǰty" ��C��JA]�c��U2-����n`��_v�s���E���d���,���҇���1Z�
��Ŋ�4���_%*��K��P���D��2��+J�!O5�����'��B�Ɗ��=Ǧq�\��<V@1	����k۹�2��3��*]x�w"q��7�f��Ӣ�X�f����T��R�)q�5SS�=���Ɏu��sU(�X�}�.��=j46;P��T�����v��H!��K�(��<JS0b���^��?�Ke�V�f���z �x�ѫW���1y��J(���O��oN(`#��UL��s7���S2�eԆb)A�Ƀ�L��Jz#�iQb,Q����v3?������']"�Ǉ4dCP#����hMx�؉h��Fz��������4{�O�mT�#���U�y!4�.[]NX�w�s4����_Qd���#����_�V)*�&�5����5"A&j,t�B�XX+��%�	\J�dǄ7L^)ˬ�謪=�^>Ľ��n��GF8[;��(g�Y��[��5�l��e���8xrs�.N���,��s�	�=h5
�e[�o@�jL#j�$40Ő�,p>�+(K��]1�f�c�Ϊb*�t�\3��*֖=k��,�����M�����N㖠^+c�6��}���3�Z?��`�
� uі1k�Zf"����^�s �%�3E�h
 LVSڈ'u�3V��W��+�?9�����%  ����j�NG�X�ŔK�ZvӼҟP��E��i���nW{��X������S�f�+�:)*�u��΁��4^��9`0R���m�Q�};;���M�Hhi[K��y^_�#�&�t���GY<P.��z �|`��$�خ�K5�Vo��*�?��됦��hJKD4������;��8I_���=�8�������q  $Ä���&�U�$'�c���џ�p������� *W6�
d4)��q�	�Q�+���g�S�Eg3��-
������V�d�b�[9�EA�̢��8]���5B:����%�w�����u�i�Z�ܦg�X_eX���i��,�\N0z��$������S��Z-Y��̎{5�FO�0pj���KΕ˥��~���8� Ru����-Ʌ�^s)GY��<C���.$�Pޝ3�db�Fg � Ł��lL�\���2�={��5�Y2F#`S
��>� 	���E;iޟ��|�jG��ѫ�]�I�=H;�q���X��U�5�mji/���b�����J.P��n�j��OH����s����f�t���X����~:��x�
�p����W����Ѝ���+�dr��4զ��?<�����Uk�>0�&}⮥�\�鞇�@��B�J|�M�a���*�� <��[?FN��&L�R�\?f=g�c�`����"yl�_}��,��߽ts3��戄G��I4��[AtH�C�!�YO�"m&4f��ܐ.�w�|1$�>��%6U����D3�=��<W�����"B@�������ђ���6��]��Oc�2kU%���ֲxV �z�K�@t�muؔ=L?{M�Oeugh�v�#T[�L�z<��&Zq3?�t� �ޙ��g���)E�Eщm�f;P��Y.������a�^<KAdf���%S������&�p>��R���SV�&(��c#a�� ����Qk�|>�A�~|[8m��f��Y��t��p�M~oU^d��3���Oō����>�y`R�ݪ6W�ױ_ �p�;dX_4[rh�� �> Dj�W�f���T5bm�h<��k�hS�]�ĳV` w�(�uKj���Z�T�OA�0")��e6�ǨBL����Q9�&c{�� ҅1�T�$�TuB�tS��d���Y��B�p�u�[P/��<�h��j<�G: ��}�'�ŵ<N�¼*��b=���=W��<�w���[�/���4"�������e�.��2p��K�U+�k�S�$"�]���/t�6�y�'N��6Sr>��/��u����7
��懃)3�6AKdϔ)��͔d쏟&;��ӹ��0�bP6����5nW@QE��p����]��:��D�\�?��y5:bی���㙂��`�z4�5�����t�͓�|7�?f��Σ 4��]����ɖ�l9���(xf�6EM�5����F#�sn��@�^�p�A[�4r�X�=/��{���}�\�L�)����+O������� }t�&�/lR?�F�Ƙ�Z�,�c��g̽?�Xv�ťzߩ��F!R>���U^����8D�T�8&�r�_?*����������u}L͙b��93�K9������������!/������&Աi��|�}�@�P��6�� h�F�����zV���w8r2���&�nM�3_yv���G[�XL�]��������巫�����?q���s�1a_�R�,����ɜ�m]Z�Ę�����/��'�Q�w���	�=	� �D/`�"r*t�B.���E익$�������I|L���ո���ւ����mi̆���_��u#���.y�Ͻ�����#d�P�~`�Y�8i��X;��B�X�!ԩ�XU~�	D�|�t�ѐV�7�n]�I]��7=.��΃�<q�Q<��7��K�y�=�<5���s����Y���Y89�i�|�en�����w-��%�j�={m���0����̨6�St�0�Ȣ�3�اi��c���	߯jz��/���������u���@nʓ��V�<�� 7��7��5�2��H?��3�{S���nv��r|4� 
+�����$IJ�)��+G��%�Zj����}O�"X�Ah�Ui�_�@�;��q������w��ɰ�w<r�R����]b�����öWtv+l���s2� ��®�uszxai�Ez�����9�?��zn�y:�u�Y�0��!�?��~��l៵���C�Bw���9dXHԨE��\!�|�F��>i[�Wʅ9��bn�"5BR�����S��#F���E�����%�����ѿ��e�s��,���^��/)p<�������F��sϻ�*����m��5y|�	�[V���y9=9�剈��d��<�L�}�8,��|�j����&�Nը2\v����x��>u�Ҁ���OV}jº!�j�䱌^����P5�����8(�������=A�D=q��8(E[�&����6{�˧3ǴE�}i��\4��T7�#
��3������'������4��V�����X�S��[~�#�F�G�W\O��8�0��ew�r���'��Q`""����e:2*	�g�{x��zueA�#ܺ�UCo�^S $���.�1׻1���Z�+q�U4�\���D�a-�� g�>�'��<L�5Bo(����t��~�w�e�":(�}���G�$�$��/��,�F�y��"� ?:�t��߃g��A��|,�;|�{!@uy>L���A�w�o�]�Xv��W�� #�=�Dl�<8�xD�S�� J�薢~�"���u}��89��u�l�{���"����l��􎿣H腻�bW{;9���W9۬Mrߡ.��]+�Z?Q��_�W�Ѵ� c�jn���-j5l�:ˉ�z P"�����jf4���e9dL����;���A7�ܹE���:��ä��r�EK���s/٨�s�H���ni�}I��mϰS�y,����s��W!5K店K�b��%>G)�*B�Y`E�hr$�����'��n����+9��L!�C���]|���I��y��۠��I�[\�4M�����h�Q@�pڃ���.��؀����/��,���B�#vOġ~@F�zڢ��>��/�/�]�����)���@�K��h/R�s��Nm�(�Z/#�YWc�H� �4A{�����&ıu�N����\�m
7��,>�ԥ��z*�T�Q�1��@0��I,�S2?���v��f����Ke�L�3�c�)�׈ƙ^�>�t��0�g2i�Ø`8}�3��T|l��Sj�N���tg�0�����mlTҹ��B��Nk�����D
'��Q���5q�_��:f�:���͠��sl���NRB�DF�c����
E٢�$��j��D��AY4f	Q���H�́�����H
8g�j����� Rew�2�i�E�4%6
 S�-N�&�����D�A]�fR|��S�ʔ���y+����Y�	��h���	�?Qc�uŤ%PW:1�̇�w�+����5�����q�
Qc �Z7Sc�}��_)��ˣzeUu��:�g0�^�&J���5�Ufb�<����?uQz-�2��P�Ǽ�x�6Z�޲�K�Q�X;��~v�0θ��BF̓�,���|k����	}�׭��CI]�7Ûq�������߭�;�*Ӷ�@=����s(�{.x�d.�lK�����ϙ��\08�ߟq�����g0���P,|?�*�w�u�w��}��#ݣ8J�ԇJa�X�H�3ʹ�0�=V��cfM1��e�:k�v���5�A�M�kG6�D������'�T�������T��DؖG�G�>d<�n���A�F�%N_	��AL�1�U��!'��Ϳ��N����PT=���I�G�M�P��$]��`<q������]`H	�n�9=6��ꈹ+ $�1lhY��l?�?<���y���$ڂ�4�ųw��\�bFC_*���!;b�kf���5r�x/5��>BK�#�z��&77s��t�\�antQ�܌4�I�p��F]fK�%n1��� L�<*�0D�w[8q�'���~���b)�޽��'����*��	.�i�ŭB����ca�:,KEAV���d��Y'��z�H�e�W�G%CC��\��D�P��F�V�՟�0����^<�?3��#�k
�6���mҷ��s?V%��y����0&#v�l���.A}F�ۇc��Rg/��
�1��?/��XFv�x����)Z�g�5�He�V���V=Эt���	{������m;�+� �o�Ѧ�p�2D�_�����X�E��
���:�
A���N۫i�ː�B��M����GY4;��WE�{���Jj�Kڀ���@�����v�A��׃|��L&]��w�=|gG�yLo�T_N�tK$]0q�J^D4���=t^�޸�s^@�P)<���m���5q�UV@}�!L"*� A��Y����9*vx�2W�nex�����D�K��yw��ZLAa{�r���R��5:�`�w�
A�=\zR�'�0'��\p���������DD2P�g�ӗR-��W������R�F�TS}=8��� FU%9ҲL�(��8B_��O��>{�o�j���=��8�9��[���KQ Z\�U�/C��݀SP�:-^�ShX�.+�S���f��#����Y_�A���n��:;�c"<�x���]0�D<t��i�J��؄�[v�Ӻ��JpG}�y�?�����ynmi܅[�3�[��@\x��h"./����/�#�A�e��v՛U��"m��x<N3Z��/8�A�$�E�:e.!�힗 ���|����;��US_�Nmr��+�FS2}^���-�X`q_O�S$|����K�&����yH��Ȟ��`�1갼XJ�	w~-�a�Dݍlo�����A��� �-+��pI[�X�<�ۭĳJ8�H&��O�2|<4V��w�E�G��2�â�E���r� @]9� ]�R�.✕.�q�k�S��5�;ۧ�c���R�����uk��`�Ƭ����S��Uc�-C����^T�`�`�]ɼ0r�W�/%��B�^��5~�8��G��/�Y�>�������Q���{��ם�� d�����sJ2 Jw<�g'^$��:c��PU�X�,���`Wc�-�vQt�?��i�����5�<xYɍ�G73����FòF��h����:��A`���+��9�F��e�b�C��~1�w~i(l��DT��!�	����Jr=q�;�Ѧ�ԝI9�Ц� E�R�|%<�<-��:^"�a�1Y�AǏ��ZM�p�XGU$4kVs�o���c���B2+��������'��5�-�a>Qsx�f�uqO�����t{дE8�d�m����8�7����G1"�X��4O���<u�q��9Z3JT�hd���z��Zc@N&ub'����3��a�G����'ȣ�_B�Fk�>�.)˖������\��!��E�8=ia��g"xx�l���5cld
T��t��<&�����?1�Q��r��L);��ӈn�3zh�z �[=�xC��ޱ>��O����Z-oB��`�gݖ�aڶ#B�eJ]\�>�Q��܌�໧��tS�a	A�ՠÓ��0���(Ʉ�:�7J����㥥��^'��T���4�Zтc��u�8�>��w�sOe�o�)GH��t����Dw}:�k�u`@�
l����6��Hƒഃ�d3��/�XO������E���?��:(t�]�Y�K�8F�ty�p��<��c]��J��=����hV���&0	�<�J�rki"͙#)��b8�����,����O��W`r���T�o�DkV �T:VS���=�ð8�K���7:er�:�Q{�"Ip|���5;���,�t�r��%t����U&;�%�Ο���M��j���Q]X���*�~�((^�`��i�e��R$�����{��{�U�t�ˈ�a��,{%}�ɩف-��G�h��������9"wK?�є#�2�&�N�(h�'�|���q��O�t�V�����0D��I��������Kw����Т�c�:�>���Y�<?Ve��! ^Sl���S~"��B��r*}۪���N~b%��@�[i��ig~'���ݍ!���$��&<9s�o�1�)��`��!��g[��8��`3�Z~���yQ�ZM���j�A��݈d��>�*(�����p�
�`G_�g�P�ҧ�� @o���W�p���b��]�߸D�±.��P<$s�A�=Պ��)|s�����l���B	sBa��s�$yJ�[X����*M�8#a *���y��[����6�1n',IQ�/f����z����8���>k��-
���?+ؕ8@�l#�`tBqO\Rk�C��:q��#������h�T��жȁG0�rVO�q��C�6�N��yd�f��xz���{�����r�J�T���<�6�/��n�@o:��-�X����m�3Y��>�{j�	f�жѪ!s�L$��j�B���4��[��=hJ�����:T煪}�q]�D�J�rOؿW*��p��sy�p׃`7,g����$M���?e��Sy��S_*��9/)E�*`"�Q���Zᷘ�i0��:v�-�+�*L�>�x���>0SF��rL9Z�Lm�^���J��
Ϻ���T7ҸNl��.��'�+z$ʅ���6�{�|?h� � ��$ɾ�[��+ŴD��5�X_gJ����':u���!�o��1_ǻ*��8��,�����O�.����B�UQ�	F��
����|��8���
Ұ@UH"�΁ns-3B�/�A@I�N���5�����V�0"6�` 6]K�����b&"�fz�G��~���9� c��ԾL]Zҙm����1Y�p�+��>����Q��p�v��$'yvP ��a��P�I�y�K�?NY��q<���-�-�nc� āېY��(�&�z��ڤ�f���;�G?CZC�����(!�����5߈���>)�:�P_'vÃ =���`:�)��!'ej���oҪ����jf����5y�OrS�i9��.����X�>4#;��W��a0%ͣ�%��`��x�\$��������!҆#��א˗�<���.�Ÿb���JٝNIdek�P��e�,�>�}�s �L�$
����}�$+R��-s��s,�Xq�����\7ո}A�o6j����=�&NZ4D}CF�uP�T��^�>����V&ǢT��
���X��
_%Ja��/��������1��+@�g3I��`���R-�+Imo��J�m�c��Է��̢�WG��E�q��qj��|��fʽ��O�S�)��e�/������̡ϐ�+��f�>@��ݐ[�3>��C��1����ќ��15��=�}H]����)��i�0K&e@fG\;D���~�H$��Q�)�=(E������^�+��]l�U2/�M��n�C� ئZ�|����j�U'��k�M��#�{�飖hf	^Z\ǒ�I[����F�&�İF�c�<�U!���09�����񎷘�1wv�;�J�t���"fl؁M-��L�������?�iC,5sO0n�}���Z�p�׳=A攳��=���C�u>��دi3�*@GZd[�-����X�sjY;	}����BF=��4~d%�s��)�;�1J��4�zs��<��`���':��RPG3P�Ţ�w�[d�寡�r<��f���x��e���~���=E�v\m��\+]N���7!E�$��LEP���o�4o8�Oz��IV�`>c8}�ϒ���@P�jJLв��Y�+ ���Zf��ꚽ�s�j�M��\���4AKT��rm�q����ߟ��qsM-�¨ĆN��8i�oi�
��� g_�:@7����{�J���U�D�bu9��7���	�9st��Ԩ��+cGЀ*��M��a���u������vb�����qZԂ1�q����,���o�,�d��ӥwFCMә������?*�x9�U�[ڝm�����瘳2���}u�)�#��W��n|\��	]ס �t��t|���S�'��HUTg���4�0B����]���Ji��u��w�k����D	� X*�2V3 ~����ؐX<���E��z��Z����
�4W�D���/��}��X}4
*�yP�  !��vj����z5�ޝFY� �8BH�r�O{�W���6���K��K�C�j7<c�����T.�A�
�/�u�}���_��^ͳ�Y����4M|�o��36�_I=�KVˠ���n}����2��8��3���Qq�^u��*�>Or`��T��Ȳ��ģ�Xx#���w0�'�gW<����i���z�5��/��3�/Z�o$_�N8�6��L�u�ɬ�����M^4����C/��k&��.�ÁA��lz"��O��R2g����X�) �?2/�=�<b4�Z���f`]o��FوH��le�ZL)�h�����7#:`���>���9�"@eEh^^�"�l�m�ɑ{p����t�Oq��MA�E�`<��= �����"�6z.mYrUN��Z<0�UU��x���>�6C�wP��c��U���fO�t`4&<�(�h5�ځ��1���M<D ){#Z�dX#����6W�|�oõ�@n	����@�|��C%Lrdq�:̕<�������d>a��aJlC8�@y�����U������ΔCq\^��ݢ�/J��ז	��Sɤ1��?��������-i���'��	n���2i}�lh�����z4(�;ed[x?��}�
����	=�]o�f0O�%~uYkV-�4�+lm~����y���J��OY�j#��D�( ��a��R�`�¹|ل� 5�d�������MG9i�d\��Q�!q~��DT~ܗ��o��W�U�8�.���ZTş*tf�@�&xq�s�`���"�㻇-j X�sa��X3+O��c��V�a�P>(��$.'� �h�$�c��������:ŧB��#��qՒ_�]ks�;��\��I�Q��������tO%�3�S5��3?L���کM$W�&��?���ރ�FMB�g3:���$���/,^Ӊ���.�'�^��16
՝�Z)�{pd᫱���P�A�TvW�4�d�i��Dm����������V6a�����e\�
�
�d[fw$�4]�D�xESV&���Q��U�3ߝ��{`5ܘ��(�f�e����_�b2��%�v�T��b�Õ2��7V7=E�!R�5�G�H�)����
�o?rH����!���`wK
+'��������2�ɮ�����N�o����E�m�O8��K�a�����k;W4�PK�mL���c��8B3��T6�$`��u��~H�ܤD�H��꡷���n��6j� ���ջ�yE�|�Z�E7]�3�������p�(
R�:����r�S�]&*���@�1")u���O��:�j͵���)2�v�p�B�fi�2�PbO0N��ɶ��&R��ve݃|NG�u��wܑ��B�����Z�)],�T�g��%_y���`�k�����b�����X�l�ӈ.�gL�@y!|0fت���M�:�֨��ܴ��=	�9�A�l��&6f�\/2V�2�6�O2���� �Z@�pQYm}���J�-R�� �j��[TxG��ci%9��|mK��ƴ�_)�l�2J
)���e�sH��͌�FZSЈ�B�Μ����1�5�����0��ίp�I��w�c�}a�M�1��8K���x��獪�c
ĸ�F�HȪ���)[M���C%�ψ�@g�4CH��'�A�}�D�PN[�B�FU5\�f�����,*�e�sl�XG����
eâ ���n�y9���>���P���1��ʵ*��T��莥���H�ND���|�V<�y���,ˬ����h)�Zb���jM��+z�SI���3+P����,ڂ`z�pV/��o$�%=�D�zB�3+�~�"vN
��eY|�ۤ]�뷹�*���3�UCS8i��H(���=k+������t���	=�A}RM�9�Z쐑��S�_kT���B��-�{���g�˃�#���6Lh��?0�!��+?�f��(n�صO��y{��5���t��[��%3���R"t"J�m�]mxѵr����+��!fjtC�O
ߑ�����L��]Et������;0�Ο���%�ڊ�F����ذ����\(��=;@(L�o��p�ܑ�xE�9A�S))��T��f�Nd�r�f������^84ּC�&j?���[%Zyh�:d&����B���������ơ��\�� w̿P���&�A�|�ꞏx��T�cW<9�~�4�BPQ�#)����JE�:�!k�Gޢ��l�T+k�@�z����Dͱ�S����#f�'HJ;�����M�3�5���Q�:Y�ð��6��0�Gj���4��cal(d^�I<�(N�2���K+� 1j�'	pR�ư-��	�1�n�mMS�`�i�������Ju\���8;�D;`�����DZ~��NC��
��f�OAQ������R����K�i�FL���a���	�5�C���è�wM��r�nGӮ�jdn��Āɢ�>YF?�㬋�9��ϡＲ���`Lx�Ǟ�>wv�d��M�y�,~��֣�_�rH�㸯S���ʪR��Tog� ��l�-P9��	L�0��R�=�����g�3Yt����EDs�9|������6�pod.�p\bof+��/�Έ�ei��q�j]5^;�������c�d��nG�!v�W+��|�8$�1B^i��E(٩��X~��|c�b��M��d�����.�٥�7�j�'���gc}֚Ǭq� ��N�#��ay��N��ص��:\���b�q��v��w�
η�����_aͫ %![	Q#��z'=`(�(X�[6�<���W��=��@j�LrN3Ƚ�k��tk�3��[�ԙ���cܭl��s^ũ�@��IFm8GjHd���>���9�e6���y��*<�c��fu�&��w.�71�4��ҵ��@�=xf��]3��[_,ѫĳ��4�`w֒����|��̈&���T��Q (��4�r��NA�ǔ+b����e��g���˾l��A��>٠��;�p�̹�qg9wM����I�M�S��8TGox��F�Y{��׏�',46K�?�>C�vE���v�?�:����:-���`XÑ����Ph�%��_*�����O~:��������On�7a7ȕ���,�H5�@T7ع0C��<7�7���:��̿���\�p�z �b�^L��Y�������6~4��c�(�!�LE5/��L������sXJW<дO�62��M�0@�Z�ZG�F�.#�H��!�r(P]����yP���[8.\1�_��S���h�;u���CĚ`���7vzt�N�~�~��!�.�W͜x8){h3���s���9qq���w�M��ڿ�����3@�S'�{P"蹍9X��l���ԃ��0��0Va/Rn�J9�/���r����~�j|S���}�˫0m҈e����3F���p
�nr|jW�}pМ��-=-�$a]��:��:X��M|:�%I�0�ǜM������K�7w��D����Y��.�h�+c'Mtp9���u,P�� �L��i�[�dM�_�V<�ݓ,C���D��T(HC�#�����vL�.<A�Iu��.+�`��6�~����m��6�p?:)SU2'	n��F'H�����z_�tƞ�[D<�D1�Gî�!���2��uӵ�0�c>��4���n�D��W\/�0�� (`d ��$�@�A������uq���9�/4��d=
�a)v�����(8>�e�ox)�k����`��"�e�I���6ȝ_�!	����##�����l�E�Zʔ?� A�UDk�.v�2h�sPu�"�c�I}1��~��kiޞ3��8&��V�����̀� ���۲|�⑑��)�T��#n����ߘJrg_CT;H������-���Y	�P������w�h-��lB�	6ī���m-)x�O��\L���O�l��$zb*���k��.#���z���䇇���u}2(�UHQ�u]��ıPhץ��\!Z�n�k.�Ar\f�T�=� ��Z��}t�X����k����0�⋸f�,=K�Tc|��2v�n-1���?R� C�|,9��Z�#�iӫ"�l;�A�����&�ڝ>'r�wȼ�		Kv��i���MS��}M���D|�"���#���!�^����&�~x��3����9],�-�5���wE�	)�<��]�E��#u��l
��*ܜ�bT����/_�2�Q6;�(�3W_U�:�g�y�wq��MǮ�������̷���Լ`�H�V`�����Z��>���:�i��ݰh����6ql����z�>������@���l��>�y*�_^�T�.�ٺ�vȓ�T������@��9_	�;B�N5H���h��d�_���6��2��{n��Ew�1�o���Y�'���E���.�i�3`�G� ?p�ci8��B�nT����;#'C�Q��s>�!�*@�Y&�Y]ȋHx S�]܆�c�70��Sdoh�����;n'I�4gLX�r�����.:��S3���	�<����״*4�ؾA[�i��Dts�!
��7V�zx{dx�`(B����}wv�E����V�� ۸�f�P�?-*�ʬ�0}����r�T�-_���1J��e��Z����B2)�K�����O����_PC&���${Ug�Itp����'�>�pQ�����Ofq�)r���{��Nۛ"; u�8�[� %Rp�k��f���}%�I${6����?��j��BL��%�4W�[�A�3r���rf�k�q�ۧ��8K����w�N���~H�o�@6����b������<��P%�0C����L���i����z�}E'�5�X���V�e�p�-(':�+K�l��R��]�@�am�4+H�h��N?�U�[VRgmD$��`y�s�n�0���t4�|ϔ2TЄ���	%"Z*��!~���hy�N��NË��$5s�
^dD�ff� ����g�J9��9W3� �	 )��4�&m�<��.Kq�WIJ�p5&%�L���\B��j�fj� B�Y�C0��,*�B������Jm�w<��k�F�+"��M�P/\�����bW�¢n� ָmW/eQ�9�
�@�ՙzV��F�����Q�g#�@\��֔"=0�4��G0�p��ψܨ,i�<#Q�����jƴ�v�Þf��م�������k��&�1c%�
z�ckST]�V�+C�w).������l-��`K��w����D�V�&F����d$SOOT��� ���Zg�s��&�q*q,M�p&Q5�]�/+���d��x3��7'�l;�k@^�;�����nj�b#�~T5Ko��~%j١ы�瞵;BS$Z� R�a&ue��%;z1���uQi����������!�z��h|gq,2�'7���;�q3�
z؟��Z�	����{���o'�:i����ɋ@#�N3�i����Đ�8 ݾ�ĳ�nQq<c4&���,j$N�h�j��_2ғ���'K��e�O�㟸vY�&
8�x�3�L���#�Y��PJrw.��/8��p
��v6����X�5�
Y�t�4���C����U
}��0�=��v��%�\�z!���s�����[�Y�/9i&�޳w��\U��M��3E�_��z�����*��~^q��ADb(��	zGMV�'ɡ�i�9�!��Ҷb��Ai_	�|4=�z�I�̼-��T�%�
�<V,�&��/Ȩ���P��s 8{���D�R>��׵��y�v: �Rhe�μ��T��=X�Хя�����j�E��:�����✟���2�Hޙ���U�!������v}ِ�#�r��.�LE>�@�u�Ʒw�5,a}�����ޡ�����@�g?�*���Ƅ�J�F���ƶ���o���7�� ��k�r���:ʸ�a����Ĉ~��Qз������	������2��mnP��E�Uw�4�P�3�IAU�}�8k����Aۄ��g����g.���-���X��ϫQ��e��|��ݍ��@�s���A%D�'|����q!��%f��hK�g�\��J$�?A
�ꒋ����B�Nr2��1�G�lȸ�>&�Mw�{C�݆��h����-�j����c���<n�zH�G�U�>�m�5�;9��N�i��P���)�\�������u�G �X����K��/"D���{Q�1�R�+rV���I�Zթ8Pa�6���;�ϫ�>q���O.PhFkh������c����
M�+ك�Zy~$'�]�.��kaֆW���g�4&|�������ʵW���VM��[��Vg�h��C�+@|��d��1#�2��-e~���N�TX:�歝 y� 0'Ҡ�����(�����6{׏݋r��
\M��a��@���U�\7�O���EL�Hޮ����hOV�ӖvYCڠW�g-�9��'�w���N	(]0��yhC��o�_���P,��n����e�dy@�"�}��d9n\�:���t�����o��t�E��Ɓ�����))�q�Si����&�����B�M�͉:�I�j��mz4�4+�0���SV�4=A:������;ǂ2���8r��#�bk����=RR?�_�����t���j��V[{�WǕ�]�bΔ�/�͂a�;��N4,q%��ءخ__�l�e�@�~���O��;�^�����(�7�}��L���ܪ ,dy?3������*�'%EFWd�֏xv���^�lI��GT���w����R�BU�{]֥�i޾�sW�n=-  !��T6NGi�p�� �6������S��yS+�dA��{��i���B�W��:�M���3m�!h��9��%�;�B���C��M���(&���5Q���|��Z}�#�c)��.��4�����b�>�N'�\�խ.�#�ٓc��\dkb�vZV�'lf�]��e6��j��RۻQ�Ē��g�������]Uߙ�Z��*�c�O(���W�r��+�NO����AAh��}##���T	��FSU�ϴ�.���#0�mq������
��.��&�-��8�~��3"��||��;�KMM?��,��oh�#� �D��%����7�2x�7/�a�������20/we��\����bo�b��<���	�1H,딀�)-���7��*� �n� �P��*EJk�Ɛ��og3_���3��4#"�O?S�ƞ��h�s����#4���40�()��e)���Ӑ��͔��M�Y
�>Fq���� 0E|�mI���N]Z���9�R��k?���*��V���
o�b���(v��+��?/Q�M��>N��M�����{�j�z����We��`>��rh�ծZDm]¡i�ĝM�O���܉U_�r�����Vi�����ܠ�=ْl3��$i����M��t�,�_�:��4P�.�)�I���w������r�W[�;��[Nd�� Jwt�L'���7b"�v91���b�-y��5L��^g,�;���.��cKk;� a�vG��U�J�.�x������j,*�w;�g���H��=�z5B�6_��mKM�v�#��#�y&"���g�Jݬ9���at��l��0$h�s_�R�ZB$UGX���s#��n�h����e��v���<!-vһB��*�ְ�?�A����U�7��L�B�"��U0p#�`�Iˤ�jw�m��*kR>ީv2_L]�9�HQ]���O����m���P�����8�������6�5Q��˯�.eS3g�ü���@�)i��i+�`~�H�L!:���V��O�L	;?mA�LSU����7�o�+ծ�|i�>*�X�>�4�~�[L�*���!�5N�j}C�����S�R�A�i�y��Z[_^^���h0�@�1F��W�F:&j~�A���F��,�r�HH`Z �˟A;E�:$ k�<g���3%����z�����47�Qr���ұ�w2���.PmQ�v��0�w$���'G�}��R ïJbaS��oX���1�_��[O7��x/5����|��1�+F���%��o%[b��ljJBIf�#�ze7��^s?��!�4��Δ"�%/�(����#�.
�WSR$�8ٮT�=�zl��d���,�6����n:l�Ԃ��(��K�r�e\b����z8��1k�=�^�ā2�	YoO��"�;���?�+*;H\��,������;��(�u��zD����ӏ��$#�Ć�qf��I�%��N�l�����cAݻpN2@�gp�&�qNf��cU����@:�m�LC���[��L��uQ����zB�@|���.��!kB'�A��v�����V$ҭ�_�	��7>��j[��X������oZ���3�D�����
�y��`�=���bqo�R��z��Q�+CtS2�]�t�0�����{����DeC�)[�H�yZ��-�ӕ5o��Ϗ�^5��j7�n�K���ʐM=>��U�R�T^��|<<7 S�����Gܭ\Y&n�]�_DwK���Wy�x�[�k��|l�\>���3��O�V�|����6j@1�R��I���)l9넨	,�G��P�I��J�}���r�����<z\`8f<��9�BVg�c�b�ŏ�s��A]K�xj�k��P�#b�f#�0*:Z�����*�.*se�E�$svv�Ѕ�sۛ���.��sg�<�i��P�5g�W���:`��lv9?x�6�����S�T ��FkK5���Q�Um	������)�� ������+�k�>1s[�&Q����whn��t�A��3���Y'ͪ>-X~�^S�_K���5k�2{&)]�� ٪y5w�솆!���-��_�����Sw�>y>Lt��t%Ko��L~��2�x/�>}3��ԣm�7�����v�D�Y�|�d�KgDK��-�Eï̸~@�&}���R����3X���Qʸ��ے�F�	�5வO��]��M�>EGf�Ԝ7GHԄ�I���!X������F L����@�q�*Hn�B�Tv��mGَ&"�e����!m�������>��X?�$«O)o]�,r2w���+��f��_[�^l ���V��Ժ�����6���p��(��"����i���iҧ��#:P@��hp��'\
Gf�B�VA6"V݆��j8Y�(�Tk���X���Qwlw9�<��'��#��ișN��ZtlM��A9�ZD�8u�.����<�~Gٝ�A������?`�KQA*D;���:�����C�Y��2��ׯ�l�[���>5�,o��_=ѡBD����t'�7�����kr�^p���Ȯ����w�W�KS,Y8�yxc�][��Py�p��%�M`�Ģ�K�Z�(��b�z���K@o���2���M#�K��܌���)v�ӄ�*�W�m���sW�h�\���6eSU�~x��h�#���6��b��un�jDV@ US�9|z`��U�&����?��;�X����86b�Bc�U�2�΂l���sc�%N��9lq1��P k�	���A)��oiM��kEzV�Oד�~���2���de����a��6ڝ�0N"5��[�_o��fƁ��.��[~���^�\�A�*�V����=g�����R��B� �v�18-_�NAX�K.(N"ar
	�Qf�U�^
�fi/%�r�Q�t�VX<m.�D�.�М	�CX[�*�t�,�T�*j��@/�۳�,a�V�+c Qժ{iv��ů��缣�����h�'��*dh��:em�y�8�<z�	�?��I_H�a9H�}���	Z��|ͩ�	�$��g9�_Z���i�@yV����FnhD�� �l����f��:% Lڥ䷠�?��� 6�&��0wb��hR�_@'���l��R6����B$p:�/�1�d�+z�u�������?�R7A*��Q�{�y6maß���]U����u(v񨅾0	��K�8����H� ���n[K��E��GE��;zfa��դ)˻ˍy�
���z=�c������M\����L���ܖ���VoM�8�=t��m���edՙ���;����K(��3Q��a��pH���g.�TS��}H���J��6E�}�~�;���W?��.[ґ�]��i��~����2�x�7J���)���)�w�M6$�O\ʵ��{�����ߐ��r(�D���G�Of+���x�G��.��v��P�#�P*���>ʇj )Vj���e�	�/9�d��d�vj�Ӣ�?�lF�a�%��B�2�#e�$7H�Oy�wRbD���d���G���}�n/�G�d{x��.��!Fm��_�N@"�3����ï8,��ฉ�8��Ύ�$S�c��ʃ���9�PZi�M�8��?os���u�ap0��|OU]�y��Y��R����+OX9��Bu�an5g�}��¡��eS*���0zJ�w0]1�̆��`C��iS�O>y��q�����6�Wc�A���8`>�Z�~E2�HY\�_�j�dwؑ�D�x`�hR�d�J�"X)��hV5���8'"�H�&z�<w}���KK�|Dɦh{�lc2�%���s�?1��:	+={�~ىՠS���S�@3�݂��a�{D~m]i�HE]�t��_H˭��Xk"�M��p���&#���:�1A��tX���'y�^�8g�n���7���wH��rSXF��,׵�"b��GH���_���-ئCfq�^5�b�K�&�F���s�>�zm�wۯ)�U���j���m.WV"t���:jz:��ȝ?�`�1j���`�,A=छ?�\�;d�̌�7�O��j���P(��+WӸ��*'���� �U)��e� �l:B��T�<{��A�O������W��ͱP��yb��hZw���f��ݭ�ݡ6�t�%�ۉ<jN���VSA�J��3��)�-����RQ�?�����\������K���W��q��>,�Ժ�� a�V��C0`Vg��,����7@rT[\ޞiK5խ��v���MGH�me�ccl�#̖�r?t��z�S
�	�B�p����1�6��x�,)y��y�׺����׹3�Röv�k���ƣ���y|���;�(pj����ؠw�-��6�=����wS���h(�g�r�M�ԖOLi��{��נ�V'kE�0����|,Rc����`����|���\��_��O�n�/k�Jz����w��1�p@��q����Pݘ�r�ɴ1��-�a.TE��ծ��o��4�I����X���qx���9�z̳�yן�'�]���6���`'�$�1�p��,G��[R9���-����gp�"�\}M�T����H�����>�"r�'a�Mv�dk���f�f!*Y5oq8c^r��I�I�R^��>/գ��U�B*�s0��`���n�%p~��Sdl,V��9U��4�6������_��u�N���Mx���g�[+��nhso��j�o��UZ���GWF)�����(4��z�L�Ԓ�ߚ�f�N�Y��|5'���G�+�z�Q��e/��7/ՠ�*^�z���i�Q�ɡ-�&3�'���C&}���d���2��֖�D�]D\�4�6ߘ��z�͍��ݞW�Q���g8/z�Ρ�I�U�Hn8D8��6��S��k��עA0�!=�D�����L�y����"��]]v8��e�kr�=��w	JL���E�*	�b�h`@6�?�+�ȝ�0��5�ğN���YQ~e��T�DjvE��-=�L@�L>C��;I�ו;U�Y�'�i "���z�/�_̃�ڬ=���J<\!��yrv�Q_�D�AQcD'���,³����e�5������/���l.�Ճ�g�]Eq�$�~����g')W�e��xŽ��#ʎf����j����bfl�&����2�S0\����v�;c����'򕻏����V�����pM����0f���a��Q�z��@�=�1��r""�zuu�m��n٪�a��J�1�lx�iy���\���i���f���b�E��f�+��2�?R����8��+���笴>��n�_��և����������������vݍ�H/l�4A��	_�az�}�SK������#��r���UpF8���j��[-_/�(��lM��J��D���b*H�Z����ɪD�=�^C�N�9�sV�G����ԫߍ΍�f�7w�pq��������q�ȧ��l����`���o��[������C��k���Erq`7��r�:ȷ�z?�NZ�L{����B�ݔ�򩼊������۵�`ڠ���xz�a�V�R25uNԃĉj��i��C�9�l�+~Ȼ�>��V���S1���-s!�{W֚d�ᚱ��j�=(�9\��3�Yk�
#o���Wo#��;����(�̯�n�4�?[�k�O�h�l��<�2|,
WF�B�<�ZE��pC_uR�]ތ��j��EK>"m�>�r���6[��bHf)ݭS�b��b���e�Y�Ǭ�oH�d��w�d�l�Y�hdx�|�rK~o	o/B��}Bu?�]5ߒ�vwx�N3��6bL��r0���V���#�%��NN�0��+� D�^]��1X��;�-Z	b�,~�����W���t;�F�A�G���- �*3��&w)��_�� �VX��}�|P�0�N��G ���u`k��)!i�{U��������6{	�C���5ƽa�%]'k�Zߥ�u��B��a
��;�*�I�O�)U��L*gS6Mt%[����
�=����2Ey�N�ر9p��cnz������t���Z���څ��N�{1`����
72Vݲ1�2��=��[�F�ɖ�������:!�*D��ѱ���{�ڦd����pm���h+��|F�|8�Di�Kx�v.�-S��Q�P��&���Z��=�@�=h�Z,(݄�X����*z��]Q�����'���b5pJ����ﯜb $*s�W����I�f&�lʫ�7��x�%�9�����h:Z�~ۏ���u��#L�Q�K	�U	��HT�Ӊؓ���ψ[ܒ{½��h�-dL??}T���,�"�r����(^��]����u*�c��V^<��XZ�o�����f��{�pC9!��BJ�e���빨n"4��`L��.��x�Agh�/)�pr�=(CI���%�*��f�PYr�p60P��ݪ�m��-��?f6x�� �&���p����(�Mzx�B�?��|v����Ҧ�ܩ�Ď����5"�~#D@F[i�S�j�n�ٔbW�Pؼ�y����;�$g�k�S�&�[��92�8[����P'�@�RC~�<�~��;��K�3�-�t5e����,����M�]5y�'���er��ˋ-;����B��ξ�'3����|��K�ӏ�	�cgțJ��u�x�q�X�m���Q���:-���N��gSt�y��-*ѧ����d&��LK�M�'��"������㗈X��&9�"�uz6���m���_�����'T� +j`�eS} �r�D�A*_�#��k�#fږ ���:�p��|�#�=���w�@���*�V�)��ϒ?����nn/3�CL6�Kn��)�����L������<�e�=�& �F���BxQg��v�͇b{IH���f�Ub�pbt��I�Ɗ�'�d.�Ę3�46�`��k�2jqC�������eN�M���w�4�9��W�bE��ӨP�׷Qg�ܵ�*��5�Q�h�X�;K��"��Ҿ{7eC>�M��:�߫���L��̮7���K����H*�C ��Q��"(*�e�� �vH�^�JNII]?&�q-�`N�h4������!���Q	X�ʁ�fa"ϣ���b#S���2�G[�Ş5S�>w�G`�Fޕ�oUV�]�Ku�q��s�A"X)O��z>�B���.,�EG�pn.��򗗣{��/H�� ������7�A'�/gBm�ʘ��ݺ���,��|�Ҧq�nכ!Uzf+���V�岘ݧ�[��A�a����o,􀬶v��X ��p!������{{��G�"�dNI�e`��L-���/��C8X\�\v����}3Շ<��;�
'�5�W�YX��V����� &kX�h��5mಱ�{o��>��lZ5�hC�8(w�I@��݄0�uM�\.<�n7����3�~�qe�!����Mƾ��~24����!ӧ��hk����.�A�9�(� M�/;xk�ރu�)�F�տ�8��d��i�,Y���M�ѝ�����T�J�Yx��·D�#�(����~@��A:��4%&g]Wگ�O�\c{�yX����� Q.}��[ưB`��DKu�:,X+o�<�����B �9r/������2	��K��YA�����&��2gՊ�"K�������<t}
��d@e�"�U1ْ�k�c�������V�;A��iW��#ϻz
��Ƃe�A�i�Z��)�ՃP!kt������>1�0�Ȳ����Kcj�NS�ӄ����ˆҊ,c�ps$�q�*�퀔Lg�֜`��xGb�͎./��`l\3�]��@��8��}x�Ȭ�A�fԉ>⪛?Y^�6�0�<'��
��ҕe�`󱱳�~'�.`+2|LL��`aX^b֡@L�h�}\[A��=��<nQ�?jb�vv�����Bu�<��t�����_�!mrkݢ���	����G{��hI�/� ���!ێЦf�OT­�z�#����C!+�_h���2���� XFz�]	�Ɲg{����ً�8Ms�i=Vr���1�&�W�����ǖ�G��q�Q�ȭp�I<
 �ޕ-�:7#kY�Ոy20C�D|�s�����+�QB+�"���$��H�H��� ؁Y�5�(O1�ގK�,�χZ�e�&ݮ큩kd�Ҕ��BeG��{��?�^�$L��������̆�ĘyJ�s~때/*sŊ����W������ln��������~NL�#���h�I�V��O]g[�sa�b�(���<L-q�]�6�͹�U����]��i�>��W��I����r:��ZY�D�, ����.����/b��im /-��8u�K��hm�j@���d@�%1	�G�����$p+/ ��n/"���< ��U�ܯnH�[�j��!�q�����3Ye	���9y����~�>��c��G�B
���|��4!9_F)��!\FUƺm
h�; iTB�F��a��#�op���|�ϥ.z���(?�8��9�c8�J�Wv��}��Ne+g�ַ���S�Kt�Q �r�qj������C���(�z��}��R{��!n�����cpZr�:<�uCedU��Z��*PU5�G�i�y*U}�l�B=mV.�D��р���g���H�vTy�3�Q����nK���r#	�r��t��sonӫ��<7��km�]�]e��@/�.������)��<e���Tq��i4���qG����G�o�L_(@�ǔ����{oΩȢ�?��h���ڮ?��akn8��7p]��T�V��F��j�z�X�.�􊁇Z��(��P3B�3�������Ď^��w�bN=����b������nLR��c�����G��|U?(m{�i<J� 7��?a�8t���*�_����������M��٣�E#F�y1����ҽo��`�W^��~�q�ͽ]�!�F���4:g\�{��Cͻl?�9(71ά\B��.����w��@1֧eO��	�!ۑ�f�S��(��7��p~��->:a7ׄ���������+���-�N�b�I��4�-Mֻm֘o/�:=cf��9���"uq,R�d����g��0��vi;V�]jҮ�|���q�����^�Ke�X���a��R�� K�ٴ{���qӗ�}q�nޗ[��$��;���˶ߑY�
�H��Eռ���h R5!53L���I;HQ�q���*7��<�B{�%F��mP��9	�� ���g�V���i0b��gW,׹��\�V�%��o���zõ��7�u}N�����YO���Pڟ5Ne��.���y"�a�^���K�%��Ǽ_s4��eF�����x'$�Z� `L��L�a�@���哰b���0�4B&�\q� ����Xl����NH~�|P؍9>�c/c�\�WlU�8+�Y)[;�/�d�J9+Pp�Pt�(��]�)^)L�͡m� u�݁�9D	��R���[�|W.�*��D��N���6��[i%��.����^����7*�E��|l�� g+�me��-P����B��˝�N��+��U-��T����g{�;l���)�����V�ϯ��G��,qX�l���~:�+�s�V!ox�~RBގ{��Z+;J��%�*��i]�ُ�>8��_nM� g)�ąX?��������J&]����j�Դ���f�Rb$�g�D8�,���%���4m���v&��3����h�^)*Lی9F�"������r� H���㰼��G��.�81������k|io~Ҕ�����	��NHA|m�X�'�.a)b:���]<�:e��G1�U���="��S����y�#�f'�@�=0;��8�@���E���/=�bP��S�*��d�ր�J˔�
ųP��6ǉ�CoWT#u_X���gm�5�]{5�Lq�I��Sfl!ؿ�I�[����������,նC�;L-9�5�c���L]eC6��T@Ľ�B� ��6R�����i@Gu;��Z�|v���\Hq��c���ڟ:��7�(�����;��+�� ��A��.ή]����=�%�|hO%omC<:�e�~e��>3<ǡWo/bh������1��;��1:�Y*dQ!!���a�?���2c��̤G ���&ƈO�˲)^�L<���e�_?��Փ���:��y�������?aR���	�gп�ګ��ܧb��mۅ(Sڶv�0*���#F�z|:#*a�2�ԟ�����u�./����&Ԋ�Kg�c$c���o.8x��@U���G]���L\�7�� �nJ�x7���e��m//�|��$�	�g�	���xS5���B<�B��?K֔q��#��F�?���Tzs���Y��a[�R�!Gy5Z��ѝno��6���œ0�^ �tD���>/̰�A��`+�K�߻x��!�j�A)hw�Im�!SM�4�]�%" ��h����sF*�(����<,�@�&�4=��N�^�^�1�Y..���@[�!y��۵61X�_�
����T���c�*3Kё�2�R�J��߫_)��<Q���@Pj<w�����X�ޖƝ�I��2���7����cy�p��'������oX��wʞ�'`�9J�~��ߌ�ov�/K�!kqz@Ӿ�K��j��!��W�}-���0Kp����W�ٴ	/���p7p~�<s�{���@�3�&`�s}s��P�p*��M@��c�����͠�|�0���e/�}.����L���z,E��/�3��SX�%T�<������
�V�\8�����,�	��m����u$~W��s����Ԍ|�����3
��Gs�d%0O��ٷD�$X��_�)���KnU����6�J� t�C�5oK���x!Ѯ�ݩ{Ϸ� ;|7�����J5��'ɟ,���Td+$ �6J���=�h� �1:8�����4�Z�?D�i��69�7��"�C�/TR;�W�[[WGHj�f�ȭ���Ѓ4���_�[��N-aޗ3�Tt�E�4�����*����<�ܡ떧�	�E�������<f��SL���%8��܃��xS�!��]K�ʰ�CI�*)��e�o/�*Ba;�W������QY��x��-���0o�{}�bI}y5/�}��QO��i;ͧ����WqO"�6��$1���+�Ћ�(�]��c��zQq�bh�D�����q����.�4ɮF���L�#Yq����qk����@�#I�d399/�Z��TF3��i	��3�����_ξw��]�즸S�R�fIpT�i�F���"��4��ρK  �BˈX;�䀅5d*���1���8P���#�h��d���T:� �W
�3��7�W��a�y���U ]&r�݄|�5�d�=#玬҃B��Զ�j+|��ܳ2Wk��
��+�_��i�?pid{�Ԓ�؊�L�=�]��X�m�Q*��_�d����g>7�G����8i�v�����L�1|�G�T�v�q"�t��B�B��$d!�Si�x3���H�)���͐ǳpTG+fD��5)q�Y�����9��X�^ϯ��SmU����Ι���O�NފA:�bbb݀��(��"|��Q ;:��u�V�-����.}.�_�&p֙���cdc��_��By�N5ʲ8"�)�=����v����F6ފ��qaҗ�\������r�K�ꃥ�J�Vw,�~��zn��޽��;�#��Ej��������N?`�	.ӬH�9��
�Χӎi�a�mvƙA�\��Z�3&�T��Cd�R��| \�z`YI�j6�)������|
ޒ,�ǥ��u3�#�vk��n�"��Y���rP�C�9�v;�{N�-���;p$�ߪt�jt���{�Ӆ��H�
h?S������ͨU �ɏ�td�|�׷�m6"�Z���m����`֨>pH|+6YM	�j��Mg\i"�mՄ�r�
Aw~��Fb� ��=�`:A�X>ę���\)���y�F!��j�zy�fy^:	3���+c1���&�����z�*K�6����D'�z\e�
|�\3�|2%qK��1�&M	n�H^�����u��xuӅ�l]���̟V����q�s���:mj��NT��ZC����8�g`�]C��7�w�$c������掲�h��69{�������{<eQKm��>��j}�Q��q8j��3�t;$z/Rx@M��W�W��ٹ��:'_з��ÿLq	�M���\�S��@S�&���Y,*��IXx]����@�=)m!�X6X��dIYg8I-�
/�HZ�ٙ6�)��徶^�na��:2(e1�E���At}�سZ�����yu���zB�Z�5��w`����`����N���~�N�=w2r訂�3��1�ߩ�;)���{�F�o)^ޢ�8���}=��,TOi�w����	�r����_��k��M�oS�жi��谸@� �Y%Y��"?�Cn�\�K8�Q;�}k)�&�{V�>�� ��|����D�0�>�����#�s�R��$ z+
���m�A��f�][��Ķ�˟���KO�W�m�_q]� Z��4��X�uo��M0�E�lJu���;��7�촞Ls����'8�S�#X��Zƣ���A���Y��=�����������|���xG�$�b�t��� ��ġ�*iX̯���a�>+ie��y2����Z��!_����z�>�@	I~84��>~C�?
���Oʙ�����#��ӳ/`���@J�cI��9d���2���vm;���b�y�T"�![a}�F�V�1��0,�_�w���q���cҺ|4�,@9�ݝ�d%G�mIU��_�b��"���ي�qx�9.1�셡�?����F��rB�}~�����X�� 2��I��m�T�?�����y����ָΚn�| �S7��\=��^~i�9�����H	=���ݾ�q�(����~�To��J���+�cS�r�����^�fyj�ɘ�@�|��׵(����u��� �4�5P<�[S�v��sծ�	N�B�[�C��V��9->F1e�;�Q��`C��w%�����i�(�TD m�t�����	��ۺ��T���4�e}.F�r���^�`���	6$����}�8^�����C��`�l�q����t��Qp�d��8��9��I�+��f���Y���(����5%5o�>�TU�`���e��,JB�:纲�	�1�o109^p>3#��5��C~z*��5��!%�O9W93��9�K���e� a�t_�K/�b�r�T�Aw�k�rt�	a@����L��ˎR�>���[x�J��E^��[���5h%!ʍ�L4*�9�����&'�� �o�̓7/�������nD�kG���(��\`e;�u^zh$�m+eRJ��X�5?Ao.�B�F
U��wb'�j�)G���B_c.:��vp��&��M����N�/������4�òN[퓶>�`#��0��B&�G���L�^C
����S��434�q� ����3�\b�Q�I51�����Hym��v/��+l���`��M�.�8^A)��uo�zP�M��'�.��v�d{�m�v�2Ll�(�Ș�կ9��U
e�R��*��	�`��`�C�1�,pY�b������hl)��������jOP2Y&��})�<A�ᩜ�I���ÆD#X tRny}4z6oݹ����Tw�7k�P4�F!f?�a�z�x�3QoX�Iv�֊��2Z0uC��V<�t��'�?fP�]В���}
�|���:[�$o$�N��WN���}��2ݦ���?4Q���A3�-@2aUx��p�z�Z�h���=���6���ȣ�7����qk�4F]�c��w`g[�Ir"l��?_qU��y��F������8���m<��QL7��G�M}� ���\�W�m+�j�:�R0:�)�|�_���'��uӸ��B�c@`wCQ!s����ktA^�6f"�J��l{�v���X��T;��
PŢD�1���Z/�=<���,0����>ּ����v��t�]L�=�;��/�j�EI�6�e�L��+��)��K6R)��9�x���ʿX��9��&Y��i`�{�
�����j*��"`��g4C� ���������FH5EH4.@��9���e#�3��9��"���E赣$�G�����<�⥃_�x�����F����d�"R��[,����C���: bġ�X��sO\��0��ý��%晃��S��Ǯw(�B�C��`�q�3�"a��M.W^kg��3�x���_鵔�nx-���yFN>V'�Kŭ"����fD/Z��K�r�i�J�
&�i��ph�" ,�x~�A����j���
�қ��ĳ��7��M�v�b(��<Rw��΀�����Y���L�++��.�e,d2*���e���~��,��n1z��u��D����&E������z���a(��܏4���-�{��a���H�w���ӋopV5j̗K�R���zXKX�!D\S�E-�U8��M�r��⡣���0��i��0���a{�a[;�j��r	@o^
��G�$�\U��(��~
{��yYV�q����Є~��m�3�m���?��e��Ibi�\<af_��d��M[}b�D퓏������N�X0�\��r��MW�����
�\�:�/� ~ ��eA�r�|c�53˷B��ֈ�&W��pk��Q'���O`/)��!��"�:_�u�mw��wa�!�sK�G�}�Z؈��~�iO��W?��k��I��m�$�R�1Q���5�5��$�����#_��{��`Ļ��-��>��k���\������(����]���C9*E+k��U������a���������{�v���(vg_Ў%v�h��{�D#���������ӊF�4�(�L~�(K����{����"���#���ݫ�]I�.����0�}�Z1��������'*�ΛV$�6-0_
�@�-���7�!�<�<��+�gd�	ϵ�f��A��/_U�9˜V�Ss��$��+1g�*S�x_/�D�<����d��_~��>Uk)0��C���	IZpw��(r.�^����{��s�C~M6��~��a��c_3�ԋiu���I���.��k���}?�&l�V�j7AJ�E�Ae�Y�DbO��e<�A
�@@����&�T����.��ܠ'A�EU��i�I/+w��]*��I.>\�N.��]�S aP��k2��4���q�����'_jX�\�!_���ӯq2�v��L�Rq���p����sC�'y��Ǹ�����u���_��]����F�a��9�4���f��6���m
��9?�s�6����uK���3�C"��`��?��i
b��*������y�I3<�Va6��O�'si,����K'�(�����?{(�9�2�ScOwd ��� Բ�-"���C��'�+ʒv�͌&�fQ�R�';'P�g�Z]rq#3�p������;�L� ���N^)��kfq�iA�f.�L߿FT�:��aA���p	
�� ��{}p��8�Ư�|��Y_�	q^�V���4��=�̟,]ڶ��%�����і�Q�DK`	=��"�(�~�ZH�y��}1�o���љ/���NLۉ��{����q�lvsD��!��C���0����lZ����A*�O�s\�o�d0m���������m�S���X�X�F�7�����HYǮ���ћ���_قe �5�(r��BY�WA�>��~ h|��6��0I58���xu��p��Z|n���4�[�8��a���-�/��M�
�f��cM;��@� �WCU�JQ��� �6&�'�
b�οm|�(U�����KV����Z��F��Rb�np��P�)�<I����������Y�Ma}6�&�?٪ۜʳUf���C�ir
bĴs;�-|f0xA`�֣m�.f��|��c]3h3�HRJ��hα��o����������U簕�V��� �%��ޖ��V1s/_;j{�mR+0���LG�ϴ��
�	��9LO~��58��&���HU�P���{"������.2��MS�x�%��������%�����Zk&�ݾ�u���h��b�l x�e�*2#��_�0�Cĭ�N�M�W�Jd��@�;D��k��oMr�\�5�!^�����kC��r'���x�{�� ��Mǵ��od�c������:Q<&Fإ4�Ci�^��@{�Զ�����8'k�[�������������L�w�iv���Te���&�E�9<�D�6m+�<���}��l_E��� ������{���.�:�I�#(� xr&���+�g��1�a%�6IA�js�G�H���;p�}]�P	=S9�|�U0Df�erY��Vz=����O�͢
35Dۍ�����#�Vk���N'�c���Y�� ��m�ny��D�'��u{�yh6�i��=Ƭ���iU�Im�*h���<��z˨;��Y3"���?
��2��ֆc��Z���[���V3�<�/��i� �vI��H��e8�/-��cۓ��,�\��8�ͤ��A�:,㒣t	7������>�q������㪮t�l2G���Z��W,�����ȳ��	�@j��p|��g�gxɕ�?��p��%6����r�_�My�/�Pr?=|]��He�hwZ��̴��(�f�7 ��Ķađ�yA���ݙ�H���m�S���H���b�ڟ��O��X�g��������N����Ps�>�$̈́�ߵbavpʩlx���Tb"��駪��z�G	gC��&� 	M��t�u)��T:����]T����c�tC�Dj���9V��@j�l貊G��Y�1'�z�]`�gq�*��Q:8�k�cbB�g���V�"c��F���d��^�ͻ]�B#?��'�4��v�ZL{�VF�v=M���_c���橀},�mOFk��J�l(l� o�	>�-`f. Wҫ��4K��7��XcvMm6^EG%^Lh����iV	0 Y���8����V������n�ڛk��t>��~�BK�sā�B�::{ķ�\$�F���5v^&&�1�56�9:)�.�����"���fKY�mD[���l�T��|�Tp��r��Y����-��M��S�6���2��X����Աz����h���ol��f8ӦJQEf	�I��v<h�\{#�kw��a31+�EP�\�woQ�z��F��ed��$Q�LOe#�x��[aa�.(/{W���F����**���Uq�O�+���)AD��V��'!�-�<�����Zr�m��f�m3 ��{�Eg�aY� ��휥��A�Q�X1a��9�B�Nۙ�y�s�%N�i#d�j����o$����f-�*�S�8��sM��^
��z���w�V��3�h�]�Tot?�ռ,w��Ij�.��L$�(�ȱU�,pbS���)�S?
-��kF��u�[��y�w��zGENb����*dn �$jQ��Ћ;P���e�ߗ�ܠ�B��z� 'V�%~��P�ϗ���wP,"�
��h�6�, �"�D#n-.��j�L��1��`�<���A+]��9;��}����

���h�~�f��7��3=�\�];���>:[�s�y�P�n�Cd�$���6�S��k��@*�vtW.>Y+�Dc��O���h7a ���
�כ�^Aí�+|>���O�hו�HU���ļ���QF��`'�^s
�Bm	d�0`��=uf�)��
�Òk�y֘��55��VYůD�m֟si����3zj%ED���#j/�9�Gy�x_
��	E&U��y/�|y?�I5�S+���/��� �a"���!�V݀�j�+���)���:�5o܊xH�
����W�+2�t|h��G�	�+���z6���&ĉ���#QnFM<L/�������H��t�Ob��C��\����X������
���k�'��-�;@��R}e�?ϼ=��
�_^U�`߀Hp����T5jw�.�KcQ�`W�v��pH!���K����?]S4Ƕ�C>�c[Q�N
'��tL��� Ҏj]���Đ��YQf��Vk�y����EVg��&��)��x������O�ȋ���? {;}�3F����u�^V-2�,�ά����:L�e�+�iT'cq�;\=[;סH%��s�knq�?�J�m��Bt�K��E��w� ���m�;�Lσ	��&-Ev���q� ��?�u_<�$%^݈29�.g�3ɩ���.��WI,�j�a�=��A�#*[�&I{,���1f�#�!t���dy�H�ȷO�旆a�����x�2ǩ��ᴨ����'�F~C-}�2N����5%GZ�P)|B* M���I.�n�`$�0}᛽b[������a�{$��zy���ȥf��}�B�Kޭ3��?�
%����o�/h��޸��uBX��hK��5=�OQ] ��a}��=s�7�*0L��$�n�*g��ӱ.�~n��A�sp`�`��x%ǘ�%��Y�u9 �q�s�H2��V����,Рɞ�Tp	�P�RKy����t�aʹ� �����1f'u[�ɠ'��-�� pB�/�d��L`(���y��A�"�1'�22b��2��2���z�T*�96��]rN�q}.4��xf���NP�'��%zf��ڤҔ~~�g:N��6��>�?g^h������
�,j�2��8w�ǻV ���%��U��>/�ǵ�c��|d���)�\7ש�7"��S\�po���h�6�U�����@w���&��{�t��g��i�h�2���AvD	xw�4I���L��245~&�}R�+�7�%lt�_G �XN�or1E:�бx��(~�lD���X� [�ikC*/ݠ�F��Wcjz&�A-���<�y�#Tq��e�8DW�q����w�
�:��ʳ{�����p)U�0�Tgw�6� KJ=ǃ�ne?�4��Rl�k�"�����������m �˞���$?�/��_��[_������Tؽ`w���UH���ųS�b||Cϴ�4~� �2�Y�����Zްܬ�f�w{�)���������D�+U�N�'��ihx�<y}`�IK�7F��]�#'EE?�jO��-�t�����YJ��u1��C U�x����t��O���i���u���\@���Om�t�N�@!n���gz�̔z�[� 9��FiΪq�*$~�c��b�$��RE+�|���M~M�2}�l/uQ6�ŋ�B��EG<�S�&�$�(Κ̈��ApD����Ⱥ�A��U}��	�G��G�?�Ю�I���m�-���f�8D�]'�f��l|��g�s�����/=J��T��f��h H�e:�^e7z��Y+G�2�İ����法��L��d�����NA�z|Zἱ]�vN�+gWhr�Lkb�P|L��o���n��"�cb��+�9�_^#�&؎$f�KH�����ʋ�dN|��l7�p�&�!v,�������	lk�J�#9��:�Nh��@�h;�������'\0���ﻝ�'RT��M���R��Ug�^®�;��J�ۇ1���몡���ߦ��x&<32�[$����sB����I 4_f)R@�wpRb��!
�E��0�Q;�9V,6o���V�ӑ�e��g.�J�i�����/I
]��DDG��^A���Q��N $8��K$;B��m�I
e%�:�$�A�s��FFxZ8�5܎Z�iq��~Y6�IPӝ�$�xP<Dn�V�A�O�IF� J]�c�^n������0v����Ax&=ׇ�3��/�����W�㡃��������O�6s�j�:r��ɶ)Eu��q �7Z3��|��>� �e�i wA��o<��ؼ� r�|�[2�]�\V`�s���,���q-è�og�9��lאN�ᒖx��(��A����|��b&������z�Q�V���|s�Z'N'Bܬ���I_���Um�,��Cm�[�oA2�Ő4
<p��>-���h�t�R��Ԁ"�)���Z�`%��5g	�ld�������'�t�u����#Hc]F>����ja|ˈ{Z��	�}�������2ԯ��Ն��n
7�A�4�߼.�6Q��r��bȍ,�W}�����"��:�g�w�b�17���\���l�X����씅Wf�:Q.E+my��ߙRI����w?�|����~}m���́�<�P��1��W�ѳ�#��eԌ���hK��B<-��'FF� \�7��!w���o�(3w�.����q�����o�}n\T8�^�������t�{,y�T䅃��$�Y��~Km�7
����ө7��4�M���D	˩t����r(��_��*��h{ f|�+O���0����c{e���&�"b�nDz��d�}��Av3�!���gF;<є��/�����`\H~��Ƣ+�):�_C�Yp�+�h=�ٯ�':|��Z�!�h��}[�Wa*4��'j�*S�Wl�Kb#ۉ��D"�$��ЦJ�2�N�e���M�CD�>x���b��;�v�ݵA��.jے���a 'ki ԓ�s�z꠺L��b9��)�`�YC���mzD�	c5,M���m �&�ٳ����)?I5��"^��bG��|ʲ5������G��:!ɣ�j�%.�8 (��\�����/b":Wm8RP���%,A.�����g'�6�Wh�Ri/�i�sg���P�]Q��¤ �}��qni�UPõ����@a���"�r��1�ǠFIK��79��P��M�N��~�����%|(/ȥq�zٻ��r(��JF�%���A(Ì�&�we8�`O��߱���o�Pf!!��N�_���A!&���q�e�J�[�}�H�z%|?Zpu)o5��&���h�՛�{��a:nj���9�	��^�\��W.����	ff��*���1�^���,���l��bŮ��uXRTG}��}\��PzP�?+ n��F��3��Mم++��Bԁ��m�.Tx�7t�Il��N#�>�9*õ}�=�����I�z(%��Y�	����a�b���&J�e�;�;�v�����_�] �R<�E�P�#p����Dk���Op��8k���hc�oO����_���D��~��|�Y�����$>��̗U4Y������Os���U�Ǌ�g&��TcZ>�#;_܊s ?�$�mnS��
���:cq��:��N"A$��2�N�����`��]�����-4�-��!��Џ7mQO��}ǈ�J%�#G/�FzbI�b�N��B*�gy��6�\h��~�+���\�z"��C6)��RL���&�P��\xe�lU��*)�.Ю��}�7�S7jo��jhw���Q߯��3��f�]������A�:�J���J�n��@γ��Q�:!�^x�\HB�j��f֊j��>&v�GK1m���)��^t���mlyO/ Ĺ<K��d�0�� F�}��R�]lNJ!��j�Pbo�N�r�	V1-�L�X�Ջ���S;��?o����B�7�i~~��T!%Q���R��)#3��YJ��6yZa����ښ�幡a��)����*+�~1^�q��|@}���������Z�Cߪ����\:\�L���v=arx_�(Z��2{�iRII6�F%圤�d���H��[~o�zOA![�4#T���b"�t�#�6@5�n�U�`+�S=��A�L�
���b�9<������&�k�����Q��>㲹b�vތ��cݏo*�t�K�x�:*���66�R�����+8.ƅ'�.��_��U/�KM�4]*$�5�#>qX(�m�e1/�ԑ�	X.�d���)-�#X��s�F��(7.�Jf5,��j"����C�g�}ڻ~�9O���2?��b����b�S�P��`M,Y�8ר�;fJ��;Ty�13���9�Cۙ����ۮ�V6�3�K$Zo,����a���E��Ɣo�Uw� H�1��"0.�JϘ{����E*���)���'���m��B��Lf�r�s[/���c"B��C�)���NI���J�Y	̖`ZH���#���]�4u,�Q~ո���Ar����K��2�q~�l;#�̈�r@)�1�0�Y���*�%�^��"8��A:�Lm�_gdg4�8���	.�i�A*nQ�Q�(�*3O����	J��"���Q�$�^dh��S�x[��Is�K�Rl�)<�BfC��&���lM��=��VGF���($XF�qԍw7��2������I��Z,���{��%ܧ�3K"0�`�"��f��;?V���e��;z�5� �d6� ��q*������!%|��4�����!������4)��%��]�K޻���c)�60�Qk����b�p����jF�v��9!]�!�s�J���|����s��$�%gn}.�\|�e���t��S�	�*
���u�Ӳ�eo,���<�b��K�_�4^�� ֽ��j�1��e�2Or?�k�X,>�oR{��s˩�`�B�R�c^y�B��qH�럶�P���/���w=��)#p�8�le��=_�c��ީ�ym�ag�,o�牙�)!�-PtV�l�i�m���uQ�7/��)�7Nꖼ�|ĵ��16��\H9 pA�.q���_�w�酐�^��<=b���-��eLn��?�)ӨjT�F�#6V�J�"i��6x��'(d
��n����9���K�H���40�ĵh��vtɨ��:k˸�ag8��LN����^ݧb,y��|.�s`����O�i_�p{p# ���;)���˓	��J�C����M�>GJҽ��0�{�rO+%�m�V�ѽ�2�i!N\��ir�&��u��7�`�M'��AS�[��$d ��h���<k��4N����1W���(�#$y��C��Y�|F�1�<��͚���
�Q=�$ߊ���l����u�wK��|o�WfV`Qdx��̀�Uْ�>\��.d@_c{����D�|S���X�x� ܨ�������)=䷩~��p�C+{�
ɒ����'�N�����O��-K��d=2���d\�j�ܮر˕�D�4к�QGUHW̓���C�]"e���лNw}*�ZO����ʬ� !e�������!���&
����~hͺXk=�xn}*�K�3!�o�1���_R��Ό.�t�\����"�v��X�:�d�� 7��/~�DK��r�RGB3eaR���}AV�^���>�*�-�����ǩ��� �~F��pr����Rgm)P����rt��U��S��/��{m��h��Fq���y��۴�U !����Ǎ�����Jەސ�Q�G�Q���a�	~��S¤M"�^��%!z0`�L{ܦ��S��+�"���s&��k?n�L!gµd3��|��K�!_�Ձ�>�������"��!G����(%��F ����Iz̊*��n�M4YH�R��
[�Y6i�韤�(S�O��{G���5tU�=,�%��b������M��e��Rb-�û���k��'��:��K����=[&�q >w<������;7���=`%��o5���D&O�nP1'nNf[��#�ϒIF+�gBا��g�gЖJ/X�۰�zn�B���sO7Xy�י�n���=<��	�[4���{@����l�H�U�n�ťo��!uH�0�x�+),|)H��@����_ �o��sQ��G�Mġ�B�:��jZ��果���Rv��/+�Z�qT�)�W��Zez���s��b�����+�Ѓ�65�X_S������1�,��=4+Qh�h�~�ON��8�Pѳ0�Ct␵|^��|�;P�FC;}z�	���l� ~��]��j��� *+/X~��������	t�>��}�NoJ���w�垕BR0�M�2��K3Z&�(u������Ǧ��3���{"N�(����6�Qۡ���s|.V6b% ��Л?��ydV�';8���k��؃�u�5�*ו�H������+����~7j	{�^�3�v����[?�d�6K��W�֠�.�L&~?@�V���������o�g���,���%��G�ԋ:����R*�8��g��tf=�a$�&(�(/6���4�ӫ>���6*M�(
Ľ.�t�T6� ����$��Ow~��b���zj��kξ����)�V K 3\�0k+���N2@����J��7�B�MP�Zߤ�mk#6�:O�qL~u�Fړ�fg���
h��YW�4~w�ζD4B	���?��n�`��h�F।��FW��d�<"k���:b*���[pVe�6u�81����������P�7k��>����b�U��z^����-� ��(��u#��h��h��*`�P���Υ�&P��=��,X����v`��5�GL���|�y����*$�~�M�Z4'aSR��Q��g�����E �GR�X�m�cn���\U��=����zX���5�b2�,�:�Z� Ԃ�@!�ё��2�i��:��!�_�E~)���qj$�:�Q��z�(I7�e�+Ac�G>��!J�^=�3��e�4��n잴��sl� �	�l��;���Й�Z�I����4��b�T� �;AcEK�f��6Ӹabo�--m[����9����2`qXf/�����o��`����V��E��b�m3P�X"��](�0Hs�������|*�iUm�Ds����S΁n�#�ͫ�F��c��:O����
h�͑�{z������d�5�C؃��̑����n�`�bH/Ḇ6�%r[�K5�uO�%��(q����&S��1���p�U*��
{���dm>m�M}	M�4h��^ݮ`�gã���'}��;ռ�L�j��^뾫��Eg� �e��*g�Y;�k�����l{߳��$�)v>�-�Y�jk����l���4�����d�,�r���l�1X��)�J ;�Ыsh��ذo�e�K'��)/�'�{�j5(�oX�Y�������Wg�$�߲Z8��*@K�v�o�J��y���"4���k�EUsJ?����n�/���������c͒����[�I,&WL�
+���p.�g�NV(��6��a]������Cf�}����G�Gp%�5���� �D�]�j[� �T�e=���;�̎'����X�P��PՍf,�,�Ye�#�����9R�
ea��
�<c�X����]߄V���2�.�n@gI����M�����Z Aג��*���Ie�%;�PV2"�J�[����"�r����0 @����(`����)�f�Q��V��0��?M9�UX��D��Q�	�(`+��MI��c	l�u�H+Qn���[�F�ޑ��o�qoai�A���дym��i�.�OFԖ��d۰�� b8���Lm�~��h�VY��k͇� đv��|�$��f'E[�Ƒ&�h��ejL���D/��#��3 =�7�|��7�O�sY7Z#~VW-"��5G�-jᇝc��e�}r�ʴ׀A�:L߮R(�:0>�£||����s}S̻��Lq� ��i#�DH��� 
���?�Ώ��V*N۸��5�A0Fn��=>.�����X$�����?�������󨞫�(������?� ��O�L���
�˄���SR�b�<疣P��nkN�)x�O����(�EUҠ���N���ܼ�G�vU>c�S�U��6v/��sj�^vIh����t��N����$�BY|�C���(�ӞM�r��jJ6s�xK���Qz��81N�$e�݄�t"���*��٤�	�#�<`���L�J�;�Y's+Mǰ.��`�M���e�tLѩ�6ôvp�mL,ȝ��+Bi�';�iY��:]�k]�%�UG׿Zx#�^Vk�6�M����$ ���:�QO�^2a_ي�5)c�S?���F,�F��U�_�8�3,�'�仫�'J�o�*�D� ���F�z��6� +�g,��R4B�Վ7B���5J�p�z��Z:,��5�@'�zY���79D��ЭyF�B	���Q0�w�n��vi
S��F��KIfʳ���뿿-�� r����H�^AT��vg����(��ؖ�=�h�p�[#��7���n�S!)�i��xw��{+���۰�GW �qr�VBm�\��{��y�����w./�N� �o���_IU�E��g���Iz����+M}=R�~�T�UVw�"����H5�������W�����X�Y����W%P���f�j���.z1��ZE9��W��x�����ƨ^�8��C]1� J��N�e<\F�T�`�q�\	���M�7E\�������y2Jږ�(3x�+�u�7�H$��a�x)y�/�W:P��cM�/�7t�V�����d�ISɛ����S+����=5$�eB�W�����G����կV}tr8M��✕"���:
I��H8��x��> ǉ,F�x(��j/;��ť���\�3S�yc���`����XD˿6[�85k? ��g�^-� �� y�|�xu�f[=j�M�Y�,Av��w-_'w#�jPM�Y¹V��(�Txe�hm(��{oz�8F�
X��m"@������<gPp��p=���v��.���~�WP�v�u:�����b�;g)U^(�|��J�Fv~��_lWRO\_�5SbSpU��'��,���� ��I&^�p�e��Ds)��P��@�V�L���3:��Vz
�~-?
� ��~����U��R������p������a�↹*�5���\�x�'YM,�OR�!9.�ź�֮��!��\a?��/�X�;׺���-�3�H�z��3)΅St����Lx����^<&{�P���������uWZr��s���2k���'�mH�W��\x����+��X�/���-G��p׬�M�r~�$�I2�XLX�*��A��D����O�BR�3U�N~��� *Ct	����4׬s ��}K&��ߠ�+�Ok>�@�ӎ��);��*o�-�Uݍ��4�� w��F�jbx�
�ꉁCW�J�5�����|���E�,hx0VR�*k������-ʫ����Ȫ���� �:w�@g�wv�DzA�)�����J)|�{����1E���ݗ#r��x�O��X�
 �����<�>�8;=K�9rJ[��p���N�UM̱0�f�O*u�6(I�/���v�sixn��K�f\�w3($��;��!���65�^P��no+���+�׬h1�����^�,�59Oj���!��3$�b[�A~�{��]�h��F�@x7���o,]�~�`���L��#�r0=KQ8)��*J.�P^:LW�ԏL�/cZ� خL���r��%�q��@>0����V��҅Z˗4A��"����3�Tϔ�~�>�#�yߌ��G
�D/����U+�7^���nxε�BeQ�J�U�r�}y����'c����=% jm��Xң�Q@l�R��rh�q�`s�n�ۻ*�"�X��L�i�0*�]�"�'�>�mmL�s�|Ä1��?#�q"/ؼ��z㸶pֵa{p|��:�X����;q,�؉!:9;E%x1$�k�:��d�3�}\Y�[!�w�k�]��4[���`�k��QK������⾤��~4�A�w̠�W�e�m
۷��p�#(�u&^V���#+;6i���L���G�qCA�i�q�M��p�ʏ��D4�
���KK��qs�?H�qR��a-w��Br�����3&T&��A��iuX->z��߀���(p(�RH�ZNL�����a��r���D�}Ωn`(lKU`�/b�f^Auy�j^��^
:�ǯp�e�����O����Ny��Ƚ������ĲC�P%������g�7�~F]�`n"�:4��2Og���#0�hCʑ���='�B�&���1� �(3��-VB$�2��$��T�U�ގ�4$�lO��TbUIo`!����Q�ڗ�����}�h�B㌫�hxo�Z�>��TIOZ/a	�o_×fڈ]��OHA	����-��{Oꂁ`iz�?k���윇߶�<��� oLr7R�C�9�پ-3��ՀҊ=�:���ARim�}��Ȓ���d ,����.�Z?� C��)E�'�gҮ�NԴ �W� ���x?��='�!��?>񲵆�^��M-�K'Yu��q�p~+�k��HJ��^梆RI�up>�'C�3K�M�N~��]@��T��"݈S�ר�N�R�L��������՘����umͣ9d��#1*@�8l�z+�Q�~�x�v�&ѻC�	�y�ڜ�Ŷ3G0g��!c��@�ik�"+�yN&�nN�@%��*]e�"L�d��6�CZ��v
:���շ.Qefo�b1V� a� \�ʊQ8B��(��I��	�4�je�|L�zV��h�������}�(vijc�KO�|$p�m 7�}Kq�/�|f�^�b�:�ɉL��B��z�a������W��H���drث��:dq��k��VB9��<��$!e�`
6��?{o�q1^��=����{x��w����9���U�;�_��Q�ӌε��ST�Oe��v���4�B�HAP���4��~��;�D�ߒ)�u��j��Z��� Rx5Y^�6~/�w4�76�@���}ϗá(�ɂ�od��0��R�^b�{�^�dUk˛��K z�xɎGJ�r��(Z��~�%1�*jLD�i��`���r�"BǬ;��j�dd���;��Ot�Ǜ�NG�V.}+��4��ݱޣd���c�>��&�)�h��i�G�q$��	���QSoX�����9��f	-+
C\�
M�ނ���0�Q���Ra��c*R�"R�<���n�ԺDq��a�����|Mζ|Ewrٖv��W���D�{O�"Q�#&R���ŢW>Qc	4LO��9j�ULc��R9���z����o�8�
3��&�
#�����C8nO-��n%� ϩ�"l�7.��o��w�r��\?8]>�kE�$ǒS|�	@m�'e�jN�b9�/���l��3��Řd��%=P�W"H)��.�t�̿E����pئ���Wp�iy]�����A��X�Bʴҝ�/3��.U>�qq|�F1 ��O����;&S�p��S���~��߭)'��i��aZs�D'>�ۈwє�'��h7�\6��p��ԧ�"�U��P�[�9��&f�-@��>t\Z��ZP�'8���K��GI�7̠���Ǜ�Q.�֍���s=%�7O��5'F� �^�S�T�C6j)܅B�U>mˠ���k*��c�a.ր.�9��qE����?�Ys���)�K���sL���ǆ,`��ӱZ\`�rX��3�P�.�E����ugPbxI3�&��8������V(t��*ӳ�?P�=q'l7?'��Pt\�<���W�-��V�Y�(���F0�[!����ӯ&�=l�t��	5�E�Zl�]�P�h2�@	�������c˷��٠���f¡� `����hm�Ɣ8�0wJJ�i��s�]]"�t��H�KJ�&��_�����V�/�J����'Sn.^��O�^g�|�̩��R��G[٦��Ăd��(��gܯD�|�8N<�mH��LT���rbhS�P����O0���&.�k�ͅ�iģ�<Z�h�;�U7����h:Bh���d�rY�q��'�i0E5Sl{�[�f���z�o��%���V�C`���E��9}fqZ@����$%���J�Q	�
�j׭�A���2�}a�cy�dGR:p���#Xv$��'d��ؕ���aQc
$�鸛�	0��w�_��zo�R�{��]�q��N�C�z������ѓ�yP�fm��lk�.�0l�Ӱޣ����������k� A`dU'L�h@@�ܷ����Ơ�=?��`R�Y�T?ɚO����jj�Ru������M�}�k����'�"�_��J��81Ό����=��x�֚�s��D�-�����Џy��e�.�j��dB1,��t0ҧ�_���]�GX�3|�.&G�ZM��)�%94>���K$��0���I}�}�a+��H�HP���������=�l��)�F�R^A�SlA�{�-����sck�/Z1Eg��t�n��'̄��n/�=�)n��~��j቙�Mu�ܩ��ɔe־0�����`�Wb)^�ƭ�+��XΟ:B�9���[X+����OP�{��\
KM��s]�&`?>���QJ	�,H���L�Ne�dD�<���x�G��m�*�1�K� �eчh�o������7TX���%�ŠI�{�����s �J>����b�u�hod��e���Lt�����ߗF2����'��k�>�3��~��r���oN�P�;�]�܈��%��K�|���ԔYt	��}]���qIL#,6j�!7�J�j���t˅ ?H�p� q]��Ђ�h�v��i��7	�:0�K��G�V�Ҁ�?��ǔ�`%}Ǝ	|O�O���Q
:f�2OA ŝ�h���T��7b�C�K�Λ���2ɼY�,q�n������)]�);$0�I+�e����{��[�sk����=v<c�i�2�gsK�5wn�����ߦ*�+���m���uyv��`>�>F��I:�"���A�p�{X�]N��T:Z�6$~�ʛ	���Į�z������2
'���xN�K��+v�{��)�_��7! }����V2�|�4<��%Z{�!g#��g�|P�o-�h�!�EAU
x����6�dI�A�\�9W��5�O����{��*>`��'(�'z}2y>�3�W����O��l��U�<!L�6���Y����4Y#�Z^o!���E&�M�����_�G�7Æ]�-4Ms�Ƨ\��
�ޔ0�.ӛv����9�ڍ'w���e �<$6y�����R�SR�����!(g����^����:��0��v��o�n�~�/�U-�na�݀���u��Էx*#~\���I�g"6�fH�X��U�χ�3���;M�չ�$�d?�x~w���0�;�є[w����pѡa��E���0�cqv%���"d���:��j{���ҞYn�d�(�esb��/N�=Y��F^i)���g����Y}�4s����բh#.'�ͫ�_�(LE3���h+[.��0�)���g����$��$�*�'Ŗj��ĵ�6;���"��1{�:��f�Mm h���wE����|�m��'�piuԝsI��v�<�̺��5�K&��4��\���֮��	�FmpF�OP���|T{焛o��]���i!��6�w ˏ�,.�0���ω��>k��kb�{�	P�%e��=�YB:{4���dI)L�|�J;H��ȋ{$���o-�[o�AvK%�C�F|���Eܶs;��y��i���wL�]��������It�~>I�f6Э�e�XU��v��Մ>T#X?%ү�����:�����`]�G$�iؙ�K{��-Ij\|ޑC�p٭�`8n��H��Aڵ�������c������eS ���ՠ�l=6#WX�׺�+�S�=x��ta��A�}��J�%h��~�o
���[Y�t}��9�UݑtJ��4�8�yY�;��*�}*�������(*�;� �O�nXj���b�5%�W�	1�>��س ��b*!�y իG��y�-q�����`�������̝i�|�(v��e=H��$�O�Ռ�����5`?�{���XM00�%������3��4�n���V#x��=�9E���8W���[�P�^�T��V�	WS"y��ܝ�'�����a@0�g?)�K��J��s�.�/�g�^C$8=]c�_�
�el+?%� RK:z�����1���S� u��x�֯�Pn����lz,��ӒF�h TZ���������*�l���M�����z�o4�U�p#��Y#��fuSI(���!�=��°���f��<޵�p=���(�����8����=�-�қ�^I������i{��U��6P�BZ\��05~5���P�ȣ�WMfvC����Z.�34D��ݻ�F
&��߹zi�<�P�m��c@6�8qJ՜�W��˦_�Jk�w�k��� ������I<���u7=}�~EPC�j&8���o�W����ͩ�c�.Q�uv�SP>m���!��G����5���}���������OBĺq20Ir���g:�����&q�iq�Bq!�j�F�*�����*�5e|�撼a��zľ���]�N���zx֐�F1yN�*���M�t�7>Bs���bz�m*O�djav�U���#�����#�\A�����QM{��_ե�O@C1�2��/��z�z��pl�)����<�v��-��$R׃��!�������M.I�k_Ɯ��X��:����?�C��-��J��\���$��X}�wRν�X�H�$���i4֠3��*d
'�96�tX���Z	%��Dhw1��Ɂ��7@B��ے#�[�eآE��t�%zC��5nհ2%�.q�Q������e�Qݪ6� �VkX�*�k`�~y]�N-Lv�1�
ɫ��ɛ�E�!���&d��� ��Ђ!��gѬ�t^�^���|��]WFa�J�5~�Iu���lWu�%]W=�}ĎZ�NO]�n�;���פ�=8����U�(lg�o��%ܬt�W�Id���T
�!�K���#���+9]�]d�&d���Ķ���x��>z�&5$��C��׼�D%PGQ�Q	܈�L�7��U+�7<`��\JR�Ksn?}U��S�w�<lL��"m/��/�����!Y�TB�$edyZ!�Rs?�KdL���;�����	�ȿq��*���)�Q`�����&����R����S2�.4����j~�����&��<3�)�:�ČR~��������HH�>��Ƀȗ�lT�~����EAd�Md�b/��ҹ�ə�h( \	.��6��p�[Ե��n������ڍcJ��9��c}+s����6��F�C<S���������ܕ�&UJz���,d��.�LEr0MT�Yo�d��D
�!	���Q�d�<�j�k����פ\ӹײJ�c\R��L�Q$kvx#�\�C%Z�c3j�-�u?#��ޤ����$H�a��$�n/�⨨����eN�$b��?y��K)�`����5?��x�k�O�̵9�v^L�P��l�f�Tg�J{�8~%�=�����ȓ�ʗ\lz���bP��)li�VX
���c�$h�SpJ��C����h��1����O�r������� B�H�v�<*�s-?×�"��� ���>�U��2�G³*֩PRj�K;<t��*����Y����<؁�X�^k�y����Ud�aiD��T�?@�h�]0xS��s��<3��So���H��_>��@�U�O��i.{ ���^�%�L�}���=���-��~�g�<7$�M2�* s�-�=���͉q�~i��@4O�Q�A�{X��Ss{������Hi���h-�*q�|�P[�Z�."��������]f\9����(�F�s����WG�N\A���3-m#���7����� ����M��^MGM����f�?�T��"I����)$��@�.O�!�9eY= /l����=��!�����L,���h,�3#���Y���,r�j?�N��Cq{����I�&e�X���v�^�Y���ѷ�/N��Yq[�i|Y�f����S����m�"���}�)�IS�/>��@yy���N�C'u<�6�=ˈx/�Zڷ����3CV�ڼ��fA�`��Q�	"���]�K�\wߙ L+Η���MO`���0E���ȿd����O�ɴ�v@W�z�62m�喸�:��._&D̯ ��[;7���bc��wL�񔠎����j:�F��M���*���*m��oQ�QT�݈�GSLOVc�P�i�FHzO=�P�sKo�]Y=����1�I�f��%J��:ף���&<d�߂_�u�����~���;	�e�W�}~˹�n�~P{M��)�-�n���4�Y�ڛ��4�>�	�dg4"8Y�++}-휯l�v+Jq�w�X��k�	�q�<�b�e�ʪ��z�G��	��ˠ�ϊ�ԫ/�Sݢ���ۡ�ӳ`�K!x�z�ቬ��5��W�t����IY��s��l���q�oC��d��$�sz	�ݦe��n~&� �˫��ژ`������sP���$9�����:���;�؋�SR����A����9�?����}�� ʇ�������8�J"~:N��O�	��t�������\YCc�0�/�1HKrD(�+y@����o�>"��~�aӋiݗLT0�	f'p���-���4wS�/�5��[�)�1S>\xom��U��o:��Hi#[��������k,�X<f�!�nHgr#�x"�rǩN�U���q:��Ԥeʹl#F(OJ���V-��B�� *ɔ=[�#�Vkp��"rѣ&ަ�>�P�K}"$��&�P�v�x��8��J�>$�u^��q���c� {��/�J߮'��	 �m �bRG��wx}>�l�t�[R���.z�6'W��^�3���\��eϐSB��OK����އ��ӿY"!
�0���bӯ���ݦ�8�r�Ҍ���m���V�I��;�����0,	���c���YA�A��z�3�D_m��C��8m.�P sj�Zw��wo�
�Z1,ݛ�"x�>M�~�?�S���)��WγU��\��zN��i�1챭p���y��(>���-�hn���?�]<�=F2 ⠄�}+������K�u#��:���Mj�e�w���q7sw���2����ڨe�}%>�`��Ҳw�˩/����{�M}��Yj��X�ŹD(\ 3�_�R'��˷^aU��l��jd9���@!���������9�y ���K�_*�6��/����t�)�.�a�P!��^��h�2�Sw��&,�)�#�L0��r�K�/ c�dL�K�������{�9͏��ܷ{�_h���K�*��P����w��e�-��^�6��r�d*�E�p�]z�A�Tf���I�-сnG�L~�N�٧���;D����{�$t%�l�]�f�"���wR�q#�I��;�d��f�����y_�<%H�}�BU�>����Bt�%���q�~��W��YDf���mw�U9��V��^��p����O9�j�.:��{���
 �g�	SJ��\B
�����SulGq���\�;���l�v��]�('RwEr���c��;�0t�,�d�n@ِ3*q0��6x�צ[�gsC;�$
ӼP���#�f<��ϢI�T�$k�����q6${B*�|;<M�Դ��0�����a����[�#�ZwU�T0�f�rE��$�����"�λ�*[���0v@����{�Y�`�֐*���u9U��d�_1ώ������T(F�te�{
r�,�I��?R����n�H�o�w��w#KUV�T1*H���T���?��*BՋ�����|�y&�슈���9�u%�ŷܵ��t(��R��r��f�k$2�`�G�ڈm��P�EF�&eȃ�uK��@��X�|���z�rឪK��N�{	���U��Y�
Z��8�k�uS����N�b���?�͛�WD��0mE[���4k�=���C�#ptXR5bH��G���L�/�#�$O�ks���r�l�"9��S�����Zl͐Q��7n�c����֮��{t[���DCX�|�Y����Q��/�Oj.,��/N��F�j�#��f����n��g�y����	q��/Z�n��8�5?">S�ߦ��c)P�}��H.��J�n0�Gr����C7[O���5gX�x�-f���B�J����/�����%�T)����^
��_���>ԓidgqw�7�Ac��X�+��K��!;�w�o��������c���4A~�(�w�.�� ��Z�=�\_I��*����FJ��[�	(�bpI��Y��:+��	���wpK���#q�Z���B@�̷{�1\��E���ݖ�%N��J�`�� ����X!Q	9���,��~��a�g����Yv�\�
r��*�����
m��HSv�$����97)R[��0pB]9S/�{=�C�lG��5����� �e�[�@��[�C/<V���������V˴���͓�oO���:|Y�/����^
�[�����+]��	qD�,M��%Jl�^T�#*�Y���P���ޡJџ�_D@���S{�]"�������d�}zB�j�+\+�c��V����A\�r�v78��k����J@x�{%�X�7Y3!����Tr7$�	�jU�e��(�D$o�D#����Cwp�1n�p� f�;�F�G7y�d��  ��{�5��q���Hʊ/ 7�n���;��k�]«IT��$|l
L�2\�<&=���!���T�:JI�7�j�M���@g�K��ztz�_ᖿN����<�PHl��˰�d=W�ԇ3`�@I�K� �x�,��l����r�n��ӏ]�������F~�;4y	��*=ݤ��^�u�����[������J�q��3	��%�`r�y浯j�[�m,��W(��M�D��l�7=�z�3p���
��!32��Y3~�Sz�������q�>���fVd�
��M��5(Y��)m5��}���<�9�<n[�|D����m�Na��%��DG�~9����5J�zNI��)��T�0��8)�' ���S_^ ,p���[��i|�����|�_:z��VVnw2|ex&�n?��V�69�dE�s49��.�H��UUL!p=�<�k
3r����zTDT��f}�i�A:���=�Ùxl���؈����ͅ�Y�R�̓,���w����uD� Eh��a��DT-v���$�N���8iJ���fS[�E��t��ɏ��E�7�L�5�E����)l7�{�n�E��=�-g9g�`��������Z�8:^$�<�f+��J�ᤄz��;�\��w�lgߴ"w_
mO-��l���Q�!Dw���}L\k}Ȝ��d�SĎPo��$@�+��Ԝ�7�v���|m;�%6��tK�x��5E��� =F�JU]O_k�T���������+n�ݤ܄�X����Z!�U�?��<K�B�SP��!�T��0����~�����W�j�V�b&��[��b��T��9���\�~[ѱ�S��6����P�D��Mi1���fH��*�n���pU�	��g(�r����C�n6l�($Z�a8����D[H4�q��k-j�_�ʲ!�5�}�� �쀋�~��p��L ;����c��M����c!�m���>��ĿV3FRo��K��uГ�O2̘d�~����ǒ7���< �8>5�m�p��m���+���/~��	=����l��H7]���;�p����x���FC<'歞(��1j�����|$�x�ь�ú\�C��$-��W��g٪ +���G*��O�o���d��|Ƅz-ww_L� O�{vk�Ⱦ�_���� ���lʼ�G�;+/�|M<S�>#珸ޖ��!��	�Rt�û	%i�2����ƫ�o|K�M)3�(�}��{CX�e��s)�(P ��!���FK�O��@��$#������2ߐ��p�G��l�r:��@�%�@=��R�o?���sM�T�PcA�wi\N�����e�%��Pڣ0���!��I��ARjI݄�����|u$�l��U>����}�YvG�=r�t��z�Z|��3F����c���ͻ��+lq���{5���v�T<��rn�^�E�>s���&b�и��h"�S�_a�����P�,���Ѱc{�ϩ����ux,A_�wڌ��&LN{w���Rӫ��>ФvM��C�a���w~��V�)�*��s7�q���e(�:��Vg�ubҡ�g�#G@j��"�S���}��o��飫:- �K��d��+�k#��������z=��Q�3ifjk��"�ź�?�`��/t�.��S�/�P�ߠc�V���RW}�[v|�t��w6�;���3|�;-���w {L�pk>7 �l7+E��nO�7��.�$G��Z�A?���4|ͷ%���W��ƅedL���$_�P~������v�X�]�DT�-�F�iOe�;�[������i���y�J�=���!�¨}�g� �y���^�'��i>>j �a1м���A%��G��_C^O�z�w�0�B��� 7t�#U�%��{򿼝J<�/գ ���IȠ�^���ba�d��1�EDOv�an�6S��(S�.������@6v��0{��(s���ط{�i���#J���D��9��.���O�<�B��"c�3PE[E���% R�#�ɦ
�Da�����+�].�d9m�Iæ��a^��T�;�0:i5s� ��%���S�d_-v*��<z�UC�&{�\S�.�^64�M�<Ü�>
��Pii�F�c������y��<�ㄈ���HewF1a�D���\���Ě����#WL�����j���d;~��%�u%���3�m�}�/ u�m.��ov��k�H �8��VPŕ�n�K�U�[�g��W�Ǎl��~��]W/v�/�d��=Y*�� 1��'0���X^�aS/����H_��2�s�����caAk?�(�[��X�����(-�|x[-*�����Fv����������W�WNު6��	�j��{0�bH�Vc��g���gU8� ��x�ɥ��B�9ZC[oA~����k�l)'��7���qkD?+R�F|��!/���eGv�,��$�����`1.b��F�9aGs��.d��H�S^'!��;�enq?�FC��
��#��1tsGۄpp�D��4RW�p��{�SH��$9�J1��rcJm$06l�Ѭ�W�q��z���䗣=�D���m�ֆ��e��3�(d�_�V�z�<@��F|bV�p��a��Hg�A�&ͽ�i����XB;�a���ه��j����P��2 ʱNVc�݊��� D��h��<&\�_����\�B�izj���~m-�U� �bkB��*��,%A1�t�s��,�=~0<��l�_����0� OO���~r�l��@͏GO$��@Yd���*jW)��Ȓ��=lJ�pv�Ft���攴?��l�hgd�)�p�����ɇ�p��@6���F��џ˿�CPo"�{v�=��lU˱���EL
>�z:��Y	Nr�\Q���)���F�/�0i�Apx�mPz���"�ؐ�Jh �x2���IͶQ���R��X�E2tsw��㐑i�G��c��� ������obD9T#�s�>tj��~��RI��h�7rѝ� �����'ר÷Fo�� �[L�W�/����0�g}�v�����1Z�Ŏ�u�j���n�o�x��`��PN��A�b�|� O�>�����"�����٤�(^�X+�����`E�_�����7#�ŗ��*�5X8{U��Z��*o�<���j<_�z�e菂��{��!�{3k�jsjT�ro���n�-'����q�MӲ1���KVab��$	":�H�
��R*O�Hh55��%�WD���n��l2"�+�~d����37�}F;H;�W���s��3��?8p��IR}'Pf�ќ�x���S8f,+b��Y�_.�1k�:��b���~��@��J�)j�qx/A�ŝHv^�Ha��#�j�A(��D%��+vkQL�O�R����*دC޲�m�04���s�҄;U�eE�7�B���sZP!�p�!:EM%Q�em�x����T�,�W����J�
aT{v��\ Ybh�ˁhcz�lጪx��U�ƾ��z��!$����r|���*���H�Ɋ���q
v�w�N�q;ui� �A�s�=@m��4����@~���O��o����҂#-n�$(�%��F���#Q'�0�\���v?6�V�'7�N�|���H�0����!�����ڶO��G=>&q�����|x�Ƃ`{$�nU�a��kk�)�/L�( �� �D�3��ms�Nn2��X+�
\�8b��:E>bC����Nב��o����^T�\%���|�,��yߜ���#d�V���$4�Zf\ZQ��t$��_J�\����$�V}�,v$�k�aH_���"��PϏ�P<U1�%�$��Cg�4���&;1j�U�%�
cA\F:Y�sρ*Z*�S���}�e���>��@X�m��4'�Z%��5�s�蛘����Τӳ���msj�GՋ�����V�E�n�a��i�26�bh�Ҧ��>30����O-Z���Z�+FPL�7���7P=K���h��3k�Á5z�e4 �Sn��.W����VUD}h��� �D�C؀�c�Q�_�]�a
z��n�_��+a�R�؎�M��<�|�^�w�5�F]$�j
�w3ݡ�%l�6��E	�|7>^}i�4���n��b
���G7�^ڑ͎��-��*�y1���=�+ޛ���͋Ԥ�#����������*=hnY��[}�M�%#ŝx�IjGə�/�Ɛ�&���u��=���>�v�	�e�N� í�xL��p�t��5Y���PS�����ܫ����e�Qr��y�Q�;�=]�k���r��5L�*���&�a�J��m�Z��<
Y����8�2�DIhNa=��$]���Q�r�l��z��D���P΁}�(�,[g�$�Q�7���+��pA�^�ۤ� ���ͳ��I�cJ�~@���?��	A_�AVU�X�hKq��?���&Eq�ĺ��L	�y�5�'�N�Ҝ+yǺɰ�����G�D�Y6�%�F�Q/v���m�+�kS�D�`��6����ľ�62�.��c��4^�w�q�E�L/���E�{���Y�b��~��p��,a��:�)�Ǣ�vN��{�oI�R�`�Z�\B�AЬX�|�Y8D{�|�ۥ9�:���F�ˈ�ҝ	@]~�:=�\�q�[���X
�3G�����
�1!Qw�*�������:�^4�;vm��-H=ͽ�@��ԫ��t'��S	]X5}ۨ�i bq�
w��	�#Q!G�Owp}\���ҧa�ɗ�Ym�������w��Π��mx�s�����$��`/��>醿}髊�3�� �����1ţ6�ؒt��гj
���K9�)�Q����͙#�F��%�3$��O8���V,5.�Q��_�<��c�{���C��J5;v�=�A.��$�8I'd�Fa����UF��ȡ�B�&�tl���U۳��m�|�C�7���d椄����;w_{��@� x	��O���sA�T�*T:���X"�+��8B��\B{B�������6d޳c Ŝ��:����X&�a�Zp.+��tޝ�^ȑ;�Ȩcd��x�}��S��-�[V��<ÝwQҎ�R��i]���[�6��Y7iR�z���m�?��S̝�Tx7�v�L����<:�եNS��.F�{�M1�T���eE��[N��U�ߞ�2�}�[&\�o����ep՜���ژ��i��$�R��3�D��XD���h<��Z8Q��ؔT�ԛ�h9é�ܷ���w�7�("v)���-��s���*�:�\M�D'G�XYG� �`4g�(bBq����Y��;	E��1,����F�h��;L��x�����.J&�y�enC��Ӏw� ����nuس-�4)�=����@"?qa��*��( ��j�����U�������`���'4�w⚤\����i5���Ŗ����O.;���	7�N�iiv%�w��x(*K��I�I�>C�������<g�\�d�V�q����I��ծ�f��v��z��3�C��$e�mi&.aC��F�qbb�~QU�j�*rĘ��$����I2uU]�k���+�1xuB��^c�U�ɾzm��ޛ	t�ܑc���|��j<ؓ��S���R��@K��Ž�R�K�<�x��/�B�eT�>��׵����kα5�!�C�Ӟ�������M�t�^�i����7Js��+�8!k�_�a�3$�!	f]"���Vl��{f���ۡ�t$��=�M����Tg�9���D�(%���K��t��MwO�W����8i ]%-5��m�~�K �q�%�r�b&��PK�{�ID�Ow��a�(�K	6��47���M��k8nLSI��zh-���|djNL88��4�r��V�k�3�s)�:$��j��΄�Q�0�[�鶪���CU�h���b1�Up���b�cd�$�r�_:Yk����2[h �
���+U�k��S��ڭsχV���Y�7��~9{�R�E`:8��Z�o�*�
��O�Rf.��J,�F�\Rx�m�߇\S����WHl�3���ƜN��<�%�2x �Z����_p?"	�s�)݇��1y��ԚB|��p_o��q+����������E��~��"� b��۲d�n�	,��|���v�jC'�Y�+䥦�B�pp����tA�����������z��$Sኆ��4�]q�8Y��)l�`E��#w�m���R��^ZB�o���Ь��Z\�D�잍b(�e	5K���^n�k'X��>�u��L�Rzϩ�vjI�i���%�:W�.�}�-i�l��8S�^{�R�\ZF��Y1v	�I3B�1�����1��D/�a�u�"� z�����Q��)�	t��I>�Ip��n��q˂�b�*,q��������ҝ���u�,a�kYe����c�d�lfv�UU���%�/TOH�N$�T��(E��%����Wm��;�"j� �9+l5�$�8{h��� �k��eO��O�P���6~�k�,[5�?���v2ڽ�'n"HԌ�*�Fi��3r �}�,�a3r�7ck߻)W����_8�K�q�aX��W��>�/U��d��I��0
��"}��z��P\��j�7RA:J���"��_��fʰC�9�3*d�B�B�x!��j��`{�����P�x�xj�w� !�#+��:5<r��E=X`���,
9��0��`�IjB�ˇ�����J	��+�F��Q'���i��g[�����TC1?;8�Y�C��ہ��N�
��?�$� �js)�3bЕЇ���d���;F�B�wwRY����p-<�(��P�ke#���;6���m���V�Y�"����\N�}�ħ�梩
:�O��쯼���M3H�Y;��%(.����2^��L(�7d�&���ɓ'��9)yR�&$�JBE�,� ��L�ߝ���%=A�L��|l�� ǁ�ET�{j�M8��3��tX�P�7��)����U��c�+?_��	�K�� ���	��J��іP,~r[�W�$>!Lu��1���ؐ�D��\�<i-o�a"����p��0*�)��~֒��,/^D������B�=����A��`B�+Uc�l�+�_4l��N�ݹ$ �H{/,��y�R�Dj���'-]��^��̮��Ѕָ�a�	>='��ϼ��@ض8k]��S͌�۬����Ɲ/'� !�� kh�^9F���"H��۷���J�k����N�,`�����+��!U,��8�8�������m�(0��E�o����u����x_?,�H'sv�H�ʸ�$K ڭu�mb����_��ܳ����US%�����[��~c�D8�՝���ۑDV�*]���@^�䚷�g�0Zf8<���B-�.zy�n��PLb'\aQ�@{�z��`v����ô��|lg�4��W��%ćV�u1r�UH������ r  \$M��YޡH/��ݔ:5d-����#D���s'˚�}&�Q<��J��|��Z�d��DÕ����E���&�O�v�K����4Y�_����=$�l�)Zz���*��x�lǐ������A����66�䷏�������FD����T]W}Y�������pX1g؏3U� d(xR$@ý>5fՔV;I�/Ղ)
�H9%W���uߦ���]�7$��uِ��K,<L�����(�����ޠs��������+JZ~Z�q/>Ͻl�k��ȥ�Z�ީ�׀�!�hm�	��.�<v�._��>���C�>���eRS�DZhh[��5��#��GCW83Zz���2��\���g�^vɻ7��`���_B�i���i�RY#	�l�tz����	��si��|A�ٚm���-�k��)@�����hPIn�q���x;+b����n�oG zf��Z1B�QʾY?�y��kR�����	��:��䦜IЖ.6�!��LQzގ��B4� e�mGJ4�r�ޛ^��r�<V�y޴����W�Ҩ�͡�
��T<����������9.7O�Z��?`���V{vP�F���E�̾pQ���_���ӯ�в�V=X|��y��w�@K�|����v�@�$���ۭL�����p̕��fzE���[l�ܴ�~��\�VdK�-(@����/5��\�愀I8���¯sn�Jz���\�9D_���E"��燎�sY&r+7�e꽎�=�]��I53[2ۥ�3�o:��rn��9�#���)z0�+�Ks,)_N
?]��g�js����Ft�9�G�0��jVR�H���e{��m3����t�_�\��̎�Z��d�/�t��[/��^�*���,��/��	�g����H�i�/���x��ߣ���t��Qm�X��͎%y�܊�ڿ�j.������3fe�3�B�@�8�i�f۷�x���]�G}��"�>��D�;���,��
6�)��;z$()#�?b�O��jT4�W�ӌ�DHS�/�N�U0$8y�^4�Q"�>�M_�AY.�QO`���пjTe�����w1���G���`���
�-�ݖ�/�K��Ŏ�|�[i���H�ր:�����XTl���X`�Ӯ���u��]0��S���}Kc�적Ï361�ٳ[�{���Fuv�ar�St���7˵(�x\�=ʜ���C<��h6���I�rzq�,�1x�J�C�8��nF�wm>b��'������j�5I�J��aPu�o.�)]�� �{��/Y�zt�[9�'�3����������	��+����5fB�����4e����^�����OO���K�?���tf\�`��-��`��J�LsNh���^��� �1����'�xXQ+J���c��W(����h#(N��9œZ�pr�"�Z���$H�x��σD8'�SHpi����y�V���,p'q�A�PE0�[j<��S���z� �`A� Ơ���(v���TǁFz��c|XE�u�{�.��.�#��HQz�Xӆ���0p9�s�~��hX�7F�FH�uyC���r��o���ߝ�C*ڽ�q��+Z���o�ܟ�5���`��\��f�F��X5�^��a�t�Rfn�r��j�(ɟg�`�f��j9����Z��g�	`1�WX�i��>���YjG��_�xٳ����HkT]�Ѽ9�TP��4a���}E�)�ni�ß��� Ǧ�S�$�n�<1�4�7x���h���ıA3�ܮ茈bd>�{�j��!/�|��\���~�`X� _e�p���e��h��}��js�B�Xw<� JdFռ��{k�|*[�W���0ۑ$� ��'�pT˛M-�^��0�d��x�&@Tmg�V�+/L�}
��h�P��1@�~^PO�8��\ߓ$.�3�ko9Y��d����D�:'�|U����E�bd�qe����z>�ޭ|�d�I��S7C����ʋ=����_U�l�u�E���O
��32̊f���δ�;ޚ�m�r�H�Z�����%?s�"-�J�ӹX�g�ϴ
%q�_| �XT��4&���c CQ£-4�mRNlM	�mRs>v�Y6G�E�՜@�#��^͋��0�ͤ��6"��m�����u���˥yv_PNL2̀� �����n����L\������8n��vL��s1����v8m��
�����l
�w����3�WZՄ2T,_����l<�K��hف4�'��h9�|�>�U�v?�����DKK�R� �/{ �[r?�J�2���L���s�	�dv����I,L�t�3���^����}۬)R#�j���9xhd�GwFBZ��L��I��߅�t�edײ���L���,���ޝ\^FA��G�KL.�:ֽ��,�K�����oP&�6�GXI�O�?�d.G�� �!�Wv��օp�;<�Ƃ�	,�f�QQw��#z>�B�2{�}A� <�)�d%F;^�N��[�#����y��P�┙U��� f�P$Rȹn����{,�4����=��t�Y�oRV�A�6U�#G�T���o��U���Rc��u]�M�L�_+�O(c̗�[�Aůy1~�hhx�t.q���Ya�S�p���BtU�3z�'ß��`3�����,k�s���ـ����XɆ��<K5�G���>H=��mF���u��c�X�sP�I�8�֓�&Ⱦ�0H~�U��7��ԞA�f���H�����?��e�XH'�K�;�or�[C��	z�$����;.r�;��>�&��`��R7^~M�pD&7p ;*o*��T(���J� ��He�9�z���K�IM����㳈�e��n�n���t��S�X��@Ay#፼�o����>�l�vc���'���Ow�M��!�^�����Em�u��j/b��Z�&��� B���!{Cb�S/Qߩ��c6�umdl�:z˞����ߊ� '� Vh5h	�w����d�t��hֻ�"byd���f�Ӹ�.e&��ᮈf,���L���If�"�-�Z���mZ#�>堩�I�&��)��ؓo�ir�y��v��7�ܪƅ-'��
�o��.��kP�3�p_1��<I '�u�|��.�P?	xJjG�����N��M�_-���| ��ϯ0P:�0sT��4�{��D��&zhЬ��=]������'��ǅ'���G�^��T�⫁��M=ł� >x}�2�,?�"���*���a�e�۟���"(��y%$����@���~���C?���r�ϊ����������_�(��lpȼ��.����R�{������8��P�h����猵k���F4�I�����g��z�q�W�m��[�Qk׿?�\����|�~HL�V�6�,5����-���_t�%,Я���eSã��n�MLR�l��b���ut��?jd}|�W����l5��uN,f^���?׬Tё!��·���V�V�*:���A�1Tk��@�w�ԣ#����H}�����R#��W�*��د�b�Qa��.���Q�̕p��p5WL��F�na~�Gh�~�U������O-� �&�n,يP�u�����l)XÜHER[�2,�Ft�I�<�N?A"��A�-���4sZ]��_�
(?-#�)U����?�LDUK�f���&\p%��`�|Mj��m�r�Ż��U���H������w����98�~�O���(mv�cK+�t�BCyc}���)�(�Ej9����	��nl�J}�P�5�ϴݮ�ǘ�m�W��N"�����Y���A@�ذe~�&���YM�-N;�؀�*�L���QS7G�3i�.��'�dI-����������%�� o����P��!N�,���D�l�\p��ܴ*�������k�g�"�^�T�N)vvGz�5��;2�Rpc|��_�^.�nq�d�VE��nv�(�p������c\S�_����~�ŕÄ�s���i���u�eUe�p-��������f+�`�>zG�T	�]�+�,j�����(��d�����n�3��0���_H�-���(���F
Q����@RQL������r���V�2l;@�~�H�$V0�D��1[JjQ�����i������h��/�RWws�x����eIn��Ngr{ �����y��<m��j9�yקx`D,	^�#
'lx ����a~��¡^
�����f�����ٲ+�h���ԁ��C��ʻ�����c^:*��9XD��u0Ey@�a�p�#�=�8�C2�XF�%@�<1b��ag�d#�� ]���؂ڿQ��@��-��lH��I �:g���;ʙ�'㺽���N�����Y�����
L�
���瘶(D��6�>����v������3�@��24�f��۞:��	E?��OF�\�_�Ih�Ӱ/8�x%�
g�^����K(m�A�r�ly�S~@ x�=�(��f�x+��ǆ��>A3/|o�i ����̬���[��%>����R7���>�8" 64u�g����qKhS��in�������a�hQ:J�]����*�T��MU�^(��)��ܲ��&�Ր���U�!ɠAR�yv?V7�[���` �G�L��{�]ټh��4�n��(��r/5����4	���#Gy�A���\�R)I�9��x�*k6����i�������Q������6[�r����HX��6��//����X"7�.v�u�����E8Dh8�9�|�a�o���ԧ�����n�/�v����Ț!�m��y��x���o���&��U.4�x�c>���n�<g�R�'dZ~'� n��=�ñW ݥ��M$Jp�0k�6wf_.t��ɞ�#e���a��X�X3����Y�{��͒!�w������%P*K�I�iy�ݩ��K*!���2������3@>�\��u��ט�;��%�냯��\$�Au&���>s�Q�,��G"R�Q�k����V5��^����������o!�J�JWw����&P���ͭ^�����
����1��n��ψP&�M�a"����w��X'C�6���"����cI��4�~b[n�`�ެh�&y��i��H�ܷ�!#�6W!�u���{��_'Z�{��?���I˕ZH:8:��녎yue�������bG���UT�i�R�[��~���X����`�X$�%���y�"��s�����b���T9��Wɇ������t�:�d߾{N)Π1�_�]�_�l�Dx��Q�Ee��h��?�/�G �6�ᢈ �װ�|�n������"���٫���v%E�5�@'.e����Y�(��R�Ǧ�k�����j��=^�uݬ�7ҍ�x m=���i�����P�~��<K��gT��/��v��҆�5��ջF0�����Î��1�M�r�)�F�����e.c#�A����ko���h��R�;#�~~�C��Pb�c@NBb����@��1C@�j�+D�
rۨ#�S#�T�W��1��y�#i�O��$o�����R;�#�wͮXs�F�5ǁ��>9�=�v3A0�O`��{��:T����l����M�����.�!�<+�ސEp͍x43�q����t�W?�Ѻ)���چMH��!A�sI�N�7�o��C�)�t�+��/M��O���*�g��v�V7�r[狚4�9 �b�����@�¹��,��ЦD�ƶ�a��]�IiN�լ B64�}�!ſyhP�t�9O��S�&����O�{��& �i[$�Q�K0�r�3+�t�.���	��*����B�R����]g��M�s�1��l(�����3
@�oi��Ƃ�B�p��u^���4O�XL:E)���r(�뗦U(�ʺ�B��@ &/�$�y�6c#X9����m�a�V������^�{� �$�u�)C���K�B���?�bF���"w;P���w�F��C�*�M[�`kӸ�@UI�����Lr�� _���r�{!|�vh۔�<� �"=�G�k�X�S����ty�����ԁx6���;�����Pu+]��oo-H��a��`$G���qF�5�����)0����Y��vG�x��.����w����s*�^�0�Yж���Vܽ0�*� z�.�9 <A=����S���m֪*l��6��pj_LwsY�}�C�j=��D1��n ��K|�n������T&A�"~VOG�MC�������J�7�2E2nz� 	���/����ukO�p*D��>��� ,~_5S?�귮Ō��<o�+Y��x�uY�-�z�>����t>zI��q
>v�t�̪}0���<9#ɐF/w��t��'9��D�Lᗒ� B�3�0�=U���hnty\1����� ~؏�]/[]lVUʗ��80���C34������gE�/^���;7² 6�,W�S|�UB��34ƣ�b(�7u#�4^9:7���k�_��}Ye�@��N|����)_.�,��%� �����I�1����̕o�w(���^��|�k�����8۪���>eoa:�F��`�6��T��`1�M�;ٙ
F�I1����dS����@�N�_��Rx�M%��Д��N4�oyJ7�~Fϔ1˱�h��Kv�
�����
�E1#�hg�����"������@���1� h����n����x��8�r��{z�*�^H����U�X��n(�o��i�g�G����*:�WˑO�m�3t		�8�YI+�Y*ː�`!�J���(�?��8"�	[���6H�#��e�8��f�)`dEL�Q�n��>�|��y��L+|��`�`�H�z>��j3˪��%����eLCf����#,g�W��w�6D�}B�I�#M<�=[̂�z���@�`�`�T�m���Ҡ����1nM��Z�9��"���=c�h?&��#�*��P�R��qW]�^*�9]�_��<l�;�J�Kws�ׅ���<�CT���ʂV�#�*�e��4D�	��B����2?,�;A"1c�Y�R�D�n�JӜ�s�(m��_�a�.% + ư��ӗ5���A�!�{�q���r�Zq��}!A�
�O��ː����Ƈ��Χz�Wt�_|�gg���i��S��B�ঋ�CS���|cC^�K�+��L?��>ۢ�W���w�}�U8�������"r���������o�����U��z�����1cm����	K��k �'P|锊RƎ���[V���N֏#f>K^�8���APYn��
�qU��b0����g2��J!ͧΧ	F�+#v��V"~Ҳ(J���Kt�t��/��Hv�����}R�Ə@Ӌ�#�I�pP���.��-�� ��)T� ���*p0�9�Z_\��~��6��SY 9�<��`ڹ���d)7������|��"���X'�MM��8�Ϡ03:�˨�����'V�x:�MD�%���o�F�nK���%�'�{�s���iۯ�U?@_>X;�*8�H�-q̻�BG3� ͆�3���$�ہ�}�Au��S\���wN�z>��t
U(��A�*��S�o�0sGy�J�D���u#�Ӄ���8<���H���
�s
�2#2?������q���1���*��i�8_\��oU�?�7���BO$���ɤ"\Y�R�Bō��B S�ahi���i��j��#��x��مV�W���a�GN�vʾ�5�Ƶ�+�iM��qv@�K�"4t���:�3'h����'^V-��[��VS����76�~�%s�8_g^���ֽ5���z3��r�Fj��&(��+C1y��t�U�{��4�<O�=�z��*��^�����Jt�v$���Z��0,Iƃ	<�:��z9��P
��A����(_l�\+�\��d�V���o��I��Y�m�?�����g+K��h´�)���OҒ�k/���p�6�����R	3������ IU8=#�|�Y��W���#�Z�2����<vw���/ѧ�IT�mc�؏39(������9�b����0�B���xxo�dc]�� Zİ!�ک��r �1�B=l��xs�ۊ����m��֝7� �xV�T-g�]�=�DEJ�R�O)�����fl>gƛ�N٠q ZF�}:(FbQ��fNh῅��8p@�c{l��g�_�|1cŨ�v=�Ҵ$������o����U����Q76Y	��Y�J*cS�����M�P�'����������H!V��r�����&e�״Ȣ���6n`���2��nt�([q5:�5��M���g6�!7��n��'ɭ8M�a{	A�x��u����#���%�Rx���d�q�A;Ӭe8I�������|G(�X�s�N;���:�	��N�v�����G
�N��_�s�~6�۽V��{�y�*V�]�HQ�rZ��O�OH29zǤ	�o��Ag�/e~`҄��R�]䨋ȵ�5�������#�"2P���9A�T׊�
u���pȦK9�<"��0n��&m�('L�J�(��o����`ʻ�����Z��x�C@GK����s����Noc �?�s�J� 2$ս
��������8N�I��P��;��"#�
oA�0��$�g����
��Q5��m��A,�D��6�̻�a�kd%����0�rDI�B,�	�\�Bvq����S�@��֖?���;��]��������d�� �� Y{��5�g;*�������#I,��܆n+_���eb��&5����F|;M*���!�s��i�宯�b�ĕ��"|a��2w��EƢ~�������X,=oR�eD�0ޒ��&xFj���:����dN��r,tٌF���zc�l$ݥ3ֹc]x��}U�\veQt6v��Z�]k��Ԉ.�fO�)S�E�(=��Z��}�<@�w�����x��uԜ\��O@��)ҝcb�f�eBU�VחJ���U�VA�=�kޏ;0n��i��!b閪(G� ��j�R�I�k,�Xu|�� u�6�TX	(�r�ú ]2��Z/7%�т�@#WNJ�׹3V~-��Ƶ!Fކѯ�gO��q"vue��i����ݛDy,��I�ZY��I/pq��>^��@�D����?Ĕ�K�n�5���k�:�S]��պ&y��Up\��2e��?x����pZ%���i��"��	��k�o�PQ�D6�9��A~~;�h�;]p�nA�����������@d��be�֠&����,�(�|�j.�U��g���{ޓ�``��^-gq�s����-�:^����#^�08����	��3H�n�H���� ~}-��ji.���`#�g��h0��Uw ������H��Lv�m�_J�X"�&N�Q	3�>�K,wn���a]���heJ;[7��p1�e"�B��Tg9�ϭ�4���M�� 9<g�z�����A[tp��Њ����%m8[�f*��ZO��f����H�ZbB��4Ay������N$ɢ>�br���u.������>/o���TǺ�_�;�
�]�v��/KN���;P[�$�8�l�QP�I6ż�bΩ���(�S[$V��|L�Ihf�SM}œ��o��8��Ax'��-���O�z��g����E��T	M�NC�z
�����քCs��yR�����62��Ey�C�*�cǆMu�|	؇V��Q���1�W�˺�TB�ByDв_�Vk�� qsgo��9��T�
Bg��[@�n�=�2��x+���ձ��#���$(�������z��Cf�U�arM�U_��oj/���}�k_Xǉ�,�R��@�5"5�X�yh	�,fx��#��1�.�������t��g*���\O�@���4���E�N�~����
ͨ�Ca5�D?��dD�{ �[2h��g�2��u�ˢ���������%��p�Fm=_G�3%y�cOC2v�6��@��u��]<���-��d�f�y��9GF��,G��Z�n����&�g.-��Z;�����Xf+��`b03^�륬����5�4;Pq3ְ4h��P{\���sR���l�PqĚ�$0����|��#�*���\���5���4�U4���M�W8��u���J,�ku��ʹ��"pt��|� K���ǀ��.:ڮ����]��?�lX���uO�_�;� �H����Y��k#��L˄}0,6����[��)��S�.�$�]��ߢ�����q��Z�So��8:�K�B��b��?�k5���W�EϘ'�@�2ĝ8�4��D����ƛ83U�>xbe(�2ZAn}\�GGR3߬gI��bֈ�h�[�'�Y:p���t�)&��E9��cC n���ɏ���薿�N�P��};��M$�(:]yպ�h5"��HR$��+��àϯڋU~xj�M��s2Rw�o�m(��=�9�u)m%�v����,�fX��I}��Z����➙'�~����0����5��U;-����)A�s��l"=�h��ZbR��$�a�̀|��<�����^-;y�+�K'H��
����1
�x)[�_�Y����V��Y"�TN��T�D�1���UN�T�]�ݻɿ�*�͒i���7��@i��F��P��X�U�v�����j�d��@-�L�p��L�3J^-����G�grY��i������@a�8T����C|���Y$���c�)��:����{�ħ?���nT���u&V"����M�Y��:2|b����
j��`�YH|����5#5����� �U!	��غ��>s�+��OI�0D��!l��q-���D���&S���A�x�׋���C-��Aat� �������5�C(ĳ�[]��]nX�%���98X���c(r�՜��d��{�nD��
�K��@��=*��r^�P�i;z���b�l�q�)�˴�9���7A�^9�یS��!cn�����yQ�,�b$��-fF,q�v:{6(yV�H�T]�t�鬶U�b�E����c�^|�����3&����A���L(�/t��M1�������=��|>�p�����lW��/7p�t�V�(c�e�\����h���+0w?�A��M�w� �0BR�E��QVKOn*��
[w0�?}�w�<Q�K��1���@��ͦ13X�*�J�16au@j�'8�~��
���J��Z.��ˁJ$*Q�@��M |��Z��w��}`A��&�^�"U�T%!P�� |���t=l��:�9�k{�|)?���r�4ݾ�b�����j�^�n�?��9�Tyf���?.;y�a1x��Z�G,`68�m��&��f̬1��hw�p!�½�4����b��A;p^�T����A ]M�At���bՠ.ĥ�(5}.)�EeC��_ǽF�}K�oGEV��@�{QU��8ǣ8�`s�nK�HE�$�#����P3�GȈ����4�"m�@[W�]J�CsX��snS�J\��ʬ�h�goE

N!e�wkx����9��z�Y ʎ�i�?��̢j����k2ml>2���bN���q�@}��7WD�v�ⷧI35��h�N��x|,ʫ
ou���3��^�p��߶ �>d�`me+��o��]�n��I�k��@ t�KD;��cy�w������I�J��e���p��� ���݃�B��<#����i��G*��-AJ�W�ߩ%pʏ�	��:'n-�{FK��������5Zs�׃vO��)t���F�#>���	�ϩ���󃤇�|�x�xyą�'{q2�FAD�c�O���L���a9L��|���j�9�\^��ªxr��$�ְ9�8�$v�	'm�U��n���Hk�r�a��k��lئF�6!ZbPW�B �?(�\"���X$���3.棃t�:hF����i����w����zt�s�G^�U�1�HA�WKSe���!�G�)W7�4�f'������cx��Sr?deU#��8�^Q�"l���5��`>͕d��K6�,��Z�{�UC��2��	^6������ۨu��U�IP*Î���y	7���u����]��,&������e�7���?�H�n��L-M�oD,��2i��Il.���M���P���o�&�������'fʀ[u��v/�V��ז���3��N�z�	���0�p���Ϙ��y�wŏ��,�Î��1�j���Q�MF�~
D/�t�1�:D?Q���A��i�~�=pX|Uj�TQ����_��� `����f�T��.�ѽ��ɦ眗��#�C�&�h(Fm�d�M�v��!��-����bd��y�HB�2��a���թ+(�cG�k�lI,�?M��.�m��'2C" ��ψh&�B�h���!#�03�M�g��.,�R:�1�� �A�m����Ԕ�k�K#�FT�(k��\
+���c�LR��x���gu�~��;�M����g�k��{��^5
5�����F���Tu����n_�-��D��K�����bh����ؼ��G�)c�o2�;��DX��(PtJȎ�
8��0��C'\t�s|�>�T����(@˗�d:����0b��#�;� �t��ݯz��@��+=M냟9F{��B��_���bDE&���?*��
e4옊������$�F�R���G���4JD�N�7�E�Iɾ�x�@�ܖ���sW ��M�H���3��b�_�̳��=�M����rC#z�&�A���1�Cj>S?���G�F`��#��8���O��w����-� ����>��ob�g��@�̶2�џ���i�=���bҎ~�<-;@�Q;h�^8�ȏ��Ar}�������q���5<��'A&�&����Y��`ݨ�1���s�5"�?`
�U)�b�w	+]$-Q�q��;���HT��s�o �{�kP��"�����)�H_���qv���$�-v;���rl�~3�����Y$v���2���G��OZkU�F��=��y@зR����d�CM�$#	���ݗ<�J�R��L��[�c��Y9g��h�|��+(���w�-��g��r3��9C��=�7�ъ6vo+����1e����(�.���\����.VP)�`=*�r�"�%R?v1>c��{I�c�i��@� ����i�	q�(�
��f��q������(��R���Kx���CfՐa0q�b  k7����V(�d�ʆ�Y_�&42&�(����Q�}�誴u�MZ��D�B�T �=3\��H4xT�ha�8����<���7�A�5�a��e �(�6��D�<L�6�p?�Z��Buٲ��q��3� C�mx�� �N���l��ob� �#��c���|C��+,�D/^�j�fb�T�͓����ظoIZ�%��N��Я�Y0}����l��`�>J�	��s��z��d+�ׯ�*���bj�a[�� �f�.�(�z�M�T��ƱZ���9��[�5��=��;ɬس��:
���P�~��N�?��ރB�\����qی7dD�V���;>���Y<�?C% �	�6����T�꭪�(1�l���U#��F}�YI�D!��%�y�5S+�/(.�U�Bb0�=�OF5z��=z�\�o��0������%:��V��u�&��"Ҥ��R��� -��6{CU٨��?y���<<t���b�f%6�QV�b�$@����Hl5���tm!@k�P��y�K�#��
dKtH��e|)��"X�]�R��a�#�r� �8��챸�p 8�{=���Շ���N�wTA�oa⎩����$v�
	f'Y�6l�7%�+y��g�jO#E`1�t_#�~|��tRi�j�J3U�۬�|�X��4���cFl����)*�ןKR�/���g�{�Ԃg;47i��S��[�#I���	�4e��þ��l;��v)n��oO9�8��)B%���)..]c����&�����,�M���j�%���y�G-ϸ�1���_6����y|+�n6�k��½�F���š��f�D��h�Ϡюw
{)Y��R�u�j�j͇��n#z���w1�[f#���D(�ڇM�$]�LR�S��$��3�0v�+�`sI�S��J��$S��!�:�<��r|�e׃���u� �1�;m�N�<��ԧ�.Q�EUbX��?T/z����XeJx�T�����6�W	'x�� S�w�?6 g��F�PX��$oA��8�Q������q�̰f]�)��Q��"�oR(?яP��,��S�rho=z6�M�NPi�2zr	>Mq8�;=3���:������*�;�������O�1��I����b�7�N�:3+���#�����>m��t��Sr-�5U�:$�&Tsnts�g����?� ��v򂩲[�8q�Lc}�1�΂β�mT���Ζ�}�A��>�oc���(Ӿ9�Ť�!�c}����'�!�܏h�K6���F6�������u��+���6���(���:iHSp�X1���Z�����'�"R�����']�5PR�[e��iD���rK9w�$?�w�c�,�@_«����q�xL�b���B���c�ǐ�d����/qC�c���/h���8���]�=��G��I���Bn���ڍ/�/2�-��ں���"����s�Ox�$\p��	���h]�Y��h ��z$"���g���י�w�;~,���Ss����c����i�ǿ��Z�>My%�fs�O2�+�$+D�/{�t�Ӗ�V�LZ#�^3�wxZk�����>��Rp�	ƅ��k2��Y�R��_U(�5t�oX��-��jɨ�c��a\=���㼉����:��1L���\5�U�L�%+�����cA��b�W����Ņ��	sT̴��9��9��Mh~�L��|2��[
����t<�(*�# `IKkf&n��J������R�����:��'���'�+�At!l%�eC@���ةo�ެ�h���{���☽j8Y��!�d���1���{¨7B�۲�L���%3���&�6�rP��(z�F�^HO���]�??���+�q)W,��o/�fTn��he߷�8p�1�DzL�\5��@6u�).]��c�����G��J�~��Jmc�w���.3�Y���5���������`c�g���n����x�@v�C�	^L���o��^���O�o���O��(ߗ
jI2��/>m���l��;	'��Cp�� ��jLWt�T�Q�f�߹��)�B�[�J�D�{��C�����tk��/K�)^��ݓn�4��1�K]H��-&��(�]c�)�����JL\-YFrWʏ�T�^�	�ؓ���qI�pXp_�����6��k!�n�_��8l�����xR��fD����I��<�9M� nB����NH23<S��!�D�N��tu�i�`�x���:p���6{�}�]7�?��O�H��rX�JM�py���F�Y���iu�|���)��X��䣣�ܴ�q�\v`Vf��.�5�|+\�]�^Y�
�C�>�M���� `�[ȅ�ޱ�>Qݕ{Z�N�yK��0%��������d|*�~�� ���@c|��B���I�Q ��^�w��6�ֈ�	ۮ��`!ߣ^�����6zR�Y]@R-��;�N�1/��t��>&��8{�U��$��O:^����m�[7����V���+��l�5>��R���*�z���g�XJ�����4R�K'�(s����G2JZw5�J=\fr>��Y]?�Q��@t᪬>���a���}U��ߜ�g��#����E��1���_�}g4݅Kv��O�S�����Q*}�V��~�u���D��l8����4k��N���أi�*�7�����˕j��=��`���4p�����m���c��*z�Qv�|!�P8p�r�S�Z.&g���,��m+������ *�O:�Ʋ��/K(����1D�҇�\;�LYm��'"��G&��3���ܴg��#傘%��lѺ�KD\d��n��:b�~SH�,l�Ü�}p��c��Hx�I���W���?h Ut�����q]�o�p7v�ô�O7���L���:��Z�]{����+C&gb�*�B���9�K�FOH���ヮ�PG��>.�*��	M���u�Yo�!�9l�U��	����uo�֠)5^�ZZ����Ƙ
ȕ���yu�S���2_�T��P��}��Bû9
88�-k��F�3���p���#]�������6Z����0[:�^�j�X�\"fPԍ���z)��ҝ�Í[�L�;Sb���h����:g���O�&�j�,��@��ю;<Ѕ*Ìx�g6w���؊rm�L8W;T|a��SŶF�t��w�����(�~I��o�aE�D2�o�}�&���R2��|�p�n�QY�T\�Iz̯�]�8� GD�Z��0a=���5l�aXڅ�N�F�-b�9+��hUȲ:Yg���T��I���#��*K� �f����N�{��9.Y3���cA����v�aj�y
@��INԉ�9(��1��7��ㄨ����@4z�K|��Aj��FBTY��&8�;�!�M������,�Q6��K��mQ�~^���&�ߚ��"O��\�6�7Y�#9�S�)m-ރx���8��/��;@�Ղ�ľ�Բ�X��RM�8����**c��=i�&�/�'n'6��>�D+7�^��Y���s$[����^�-�q��+tӐdY,=sM7�G�k�X
�R���/*�D��(4>6����5	:��D\�vW뷲�F��yd1�$��^���GY��!ǚj_|?�Ԟ��זd���sa���؍p(�僇�����8�崅5�c��#"�)@W3�g6��a�N�
�6�bJ�^Tض��˵"��A�3k�ڄ^�d-�����I,fwhL�7�DA�x��pcg��+�S����I�K|��b~�R �q�e��4qL(cA�6��X�*�Cu2se�?^���9/��w0��x��sq�y�)`$-���y)�La4�^�lq'�>eli͟"`9q.�����˪CC��ڂ�*���_9��y>���1xj����;@��mo7Q���w�;�
�:S�Z�߽��A�㊽E@�g�	*�����e \V�����#uuݵ�qk��4$,��'�}R#�j=��4s���htV�bXsr��	�36��&�2��g��lT?3�Q�-�@	|�=O�R���{k��f@F��?�r���p+%�^��r1ېTG�ޜ�d�~%/�}�����NC�$���+v�MdYQ�m�w���]֖3>O9�x@���R�� х�l�ڃ�ᄧqպ��s��j���r�Ʈ���}o�	��0�f|$ROK���z���@���W���W:��A1�.�c�m<W+Av`�d����+�ý�SOV��
p�TyV-�A�$�\ͯ�t�ai1��gG�ʄg��,��>���0x��F�8Rr�n,gc1��nm�86�Xɦ��=�e�bPU��(��@B.��.�u���S��_��L|&R�!��s[��X��b6�)F����!+l8����^���Mv�%s� ,v�>�r��CS_�uJH�f�<Ӫ^�V�W!�:X4��m�Ьžփ*D�2K;���p�@�WC�+��9���c��Vo��z�+�ź�Nq��m�n(��U;�<r%�ǭ�h�).�_V�{}\|R�>��q�Wd��ڞ��S�1(m�ڈc�`y�*Fϲ������ F����ar|q��B�]�L\c9�ߝ|'w�:�����i7G�<�Yxݛװ��v�	h2�S��d�L��������{y*�8����L�Z��,����uưzF �ꇱ-���%�K�)W����;]*C����пW�P�@Vδt��	^!������6��K_p�(���4ޗ�K��OV��Z*��o�{�
4�
����JY�gT�QKfK�+�b\/� ���ﰐ�)�=Š^#���5	��l��')��sت�ƔT�>ƙF�#�s���F�ٶ�Uǰs)5rD� f���h��:Tw��ʭ'Бփ!l�>Y�bz%z~�)R�C�z�g�������2��ӎd�+�~e|�CG��m�͸1�f׮�(��y�����аؙ<���qf� ��iE�����'
�RkV����VG�|�-J�$f6h{�5G�̦�%��#��q�m�X\��]��Dǐn�>�%�|��ݵo��p�y�SQ�i�{]�L�m�^Ƹ=��9b��!��"e���������y\��
#pJy�<�r�����9(�Rw�D΋���*a�'eЦ ��TJ�{�1N���E�8M��SDm�@�Yn��ٸ�:�N��'7���gA@�j�l�P�ʨ�#b1=�I�-@�������΃r�{֖� ����ӧ��v�w��C��¡�H�@.ף��R4OfK7���!Et��}l0ZQ��G]���]$l��yL������6���Ym&Gn������}����<W4;/��Ԭud	��&t2f}̨�Ǌt��(�E��D��_��BC��a�Z��߆��G'��|O<��͇pׂ=�+�d$���ֳf����a��>��@�:���K\ϫ��2(zeK�r�L���Z��T���6�}k"n^��r����
�.O��7u��!����o��ӣ�p\$ohH�}�O�GK����j�ɚ��M��Y��+@���O�TLk���!���n�e��8}��Ri��b`NjS$���`���S��u3�^,��1����zp��[���� ݁�o�+�֒>a���x�0[�r#%�D$�V+V��VLG(xg`�������/ �7���'	oj���'hK�>7 U�%���y���Z'؝��(>�gt���^�����|i����P�~���Kz�i��#y*�̓r�ɋMg;d1x�֢���şeHN<Pc�����ߐRn�^&��o�M?K�WC-T�&���H��Y������ێl�{/�T�K��2g�b*l��T���^܂D@�۞����A����`W�pe���@E��wV�|�p��ۊAL�%79j�WИ���~��@���*I|�^�mU��V�O/�9�5�d�G����i�]o�Ab[�ZsZD�ȡ�tè����XD�鱂�>K�Ș�i>�.��EO��q�u_n��x??�������'ژc%�F1d�(A.�26��7�I�
'cy��;�Ԯ�[?{[�v�ޒ�
�^��M݅����!=��V��ƢPM+S�;][t$<V:���M�4��hՑU���gY�K��E {��ͣ^�v�)�r|_S.�5X-l���fpt�#ֺZ*i�ϸ�{3��uI���bQ��A��G����Q.-ӹ%��a�7׬oɺ��ɫz���ș*�Qʄ��� �\�O*׿�E��S笥7S}�0��B+`EC䦎�v�\���f�JO�i�0���Q����h�Fy,����~��_K��4��n0g'�R;~�lÖ�wt��)4��ߦiHҖ')L۔��J� ���D�U�WT`f�{���+MEP��:�=By]�+S�Sr�����֒즁�_�^�?^�:-�ť*�M&�ϵ�N�c�@��Q�>(�s�s����ph�*$W���KQ�����g�R!��+�v�k�{焬����'\�7�<�x7�����V"�/��T�� ��]N,q��E��|4��J�R=�-u�!�O*J�~ְYB��	>�t%����}�x�PkbWt3�ؼc��Q�$�b�ME�mՅ�+�<E_|�!v|A���o!1��:�Ӫ��������|��\C���(�!��etL�T�IN!j}�M�K�Q5��J����MՄAI���U���(z~��j&�U	�\7�%�bT�5���^x��Yр�޽�L��O�L		�����V����!s��aV&�mL��N�������I�p��5��!���n��T_9���P��W��R�,��X�O�:��<�o�dL����Ӆ�� ���N�����~F��-�o HL��[�����!/�����YDB��8f��*�'>��A�q�6�,A+E�c������t[C�Xx_�n�'zhg��yӝs��Q�%At7"]��e���J<q���1�N*�u�?R����A�*NDt2&$�p�\�YġD�Z��pr[��m��m�k�DHH�𓞟݆�
������{�|`ef��z`�oΓ��æYջ��<�})���(���3D�oPO4i,X�GH3@z���?GI�p%Q-�1�=~2��&����݌Oi���JΞ}��!�Zö�!h�tWjL��씝��X i���� �ԏ7(�`rP�<j�6h�ʟ�����h*�OL�ϿvjnD�y�8f�mv0k��_/��O�|�l��� ��-?)
̕Q�Bd�f3��e�~����l��w��+<����W�I?5��4B��|ы��$"á/>WP*5L"��j�)DjWeF�9�b�`�x�"R2�%�/�� ��B��Va��T���2*GO���x�PTm��%x���[�=������Q�D~V1�dWhhz��]`�ˈ���~���*�L`�4tvu=��T�*��8}+w �Kx�j�0��vۻ
�Yգ�\��Mp)ˣܣ��@^;��'d)�u�3��̏wK��x<IRpae���#+���d���rH�f8�g�G������(,P�.UH��S/�D������ǯ �>��� )�-'� �glj����5�+ #V�cP}�#�Ot���&�në(�L�RC�
֗���=Lئr���������@юrhg˘A�Z�Qk�˴��T��Q�X��p��+�t�	� T��v�l��@���u2�����i胜��nf���1��:�s�|��yT�A��w��ZO�JN�]���lѕ�f�Q���N�1L��F����h�ᾼ rKv`��y�	t��{��^Y�~���~��F���q��C(�>���1��C�����`WeͰ���|�aU�CQ5�R�FΥ~u�G`�T�3��4!PH��X.R�a2��cU4��{`$��OF�l���"��x�l�a
�i�"�nG�"�؞�K���9xϽy�o�}�����S�"�E��a�s�aH'�Jm���B���(�龒_�Q��v����>;y��U�0�@!jՎ��E�c��j�Z�b��5.`����"U�JV��#���U}u��s�ɷ]*��&��KN��O�+T��M����4<���(���7��}�+�i4C��uZb��}$e�4h&�gQf���a���*�ၮ��ؽ�s3&�/�� \&�����3]��B�~����N\��������#xk�7���E�\G�T�](s�h��ە�G���W��*i<��p�,Tr�F�X��Am�)>C�*^8����?AsТW1}	|N�n�|�� x��F�GF/-V*OO+{��]��5Ӕ�03�972��}ՖLRbFF�=�k4:���$=^w�͊��Վ��0o�[Y��$�a�4�(�^��F8�i��!����k�^8�D�����T�|����]�.X����ԙTs���P<t{0�	�y0+�W���IF	:$\�L�I�aI��"dr���̮�h���ۺK�h<p3[�����ѯ�Pq�n�l�U/��$�!�J/����o��Cw���ro�e�`վ�ㅨ٨$a�(�X����dC;��0��^{����}s�Z�Z+Wk��TLg�s�|(a��5�d��%(,��"0� %q}o��B����|�hu ��~N�����DV�¼M�m�DhO\ߜ��h#T(U���a|j�����v*�=+���wx-����Ĭ��v$;�'��I�CI��_F��p!Wr�X�,قc���x�گG��z����b�j\������Y�֒�2�L(��پ��<*1s�?��(�3��`K$ ���r����k��� ��ľ���p�����2q��/��%3.L��5��(\K�e=Q�it�6�9'�o�<�UD���.Ȣt��ޯ��G��'���yg͈/��/�Ͻ�ιf];�#�B�ڷ�k�<b\-��i�
zU�5��bzN��!�
��}`QI^��>R�td[(���<?ʱ��nt����#<��y@�4��˞��OD�|��cf��>:욨��)��D����
�AL���TW����H�F,H�� =��J>Y�����w�)����'��U��c�Q;q'uL���z�T/� �4"����t���!�v�P-ny�kcv|m�w/"�1�*;�Z.��&(�<:����?M����t��rb����)�0½G����O�$�DR㷮H�dFu��9�i�7����������^?q���_��Ӣ��SѦL2W�Lry:�<����0����G#t�;��d9�vs�3��v�:�|��<�hv�����/KCL�"����1~���:��XeEUC"ڨ��VNd��!�ڢ��!9��I�|�2�-}�q��u�`��aU{���K�������9�U����22t�������SAf����"��Mcy��/{{
J{_�_�;J^L(�q�m�2�`ݸ�kԚ
W�*"%�7�u�j��F7�#�����l�G`p���I9��^��F�f}]��@�!�h��IEKd2n��W��������h�dao�du�X�A�-+�ƼM���;�R��!�F^�u��?�Q�yK�j)"�2�`V�z�bϽ��.�.j�򠕸͎q=|�T��t�9t���_CB�B���)����w�'YΧ{3�˄�-��_J������\���$��c_U�Ǔ�*m"��8��*���Y��u7'��C��ٹ�����s��wK�Z�/&���<[H�M;���p�j-u���ٵ	5�����!��dAع���4h�o��M�f�r��~��4_��*MN��c�AhM��T��q��wW��$��C]���S�h0�m��ev�"��G<v@8%z9E��8_���_B�l_�o��a��)L_����0�=����y�w��:2��|��n�s��6�B�8�W8�A�C������(�q��P�D`�������yC�ow�QX0�%@�j�s�3��@�%�A���iV��5�U�qR�YFy��D�������!��'e'7#��������L��-y�������%%c>��
��bQ�D/�(]�O��YA�t㽁�-���Aj��U[j�K�էnܒ��$�kC	��p���j��X�4*:�n4�mZ���z�`��0 �w�p��5�.Ћ�e���7�i�����.C��_���cr����h����pz�Bk_��{����°�I|p�Q�up=uqh��Q7�*8­^��!}Y+;���}��[�zf]N�=��sX���.��Ӆܚ���]�	�;�J�a�?���O. l��˔�;�,��:��"C��n���&���]�ib� ����	��a`}�Β�����S��ς���M�,�_�ڊ���^�����f�������3�Ne:��ة�2�q��~�S��c(���*:���j$��!���j���'8Q�s-�v�]�|�!����ȱ�`	�b
���~a-ᾏ3�fr_;�-��Y8�%H���daj`�j!aZ��[r�Q��M�E�BqR���?�;���S?q� Y��a���M�
�H2USw����,+������[m.��`X1�eD���/j,7�d����|����^���Y��ʼ�i��^c��l���J�-�?��Y ����jѡu��$2=�i��u|R�ϒ~J�& �?�<��&$�@�٣�ÔE�r '�2���S�������	�h#֓D�����������L��	A��f�<��@�w��+o{���[��]<R�z���ݦG�\5��I]K�Q֭=��7Q���$�b�e�^��|�$���1���G��$Z��Y.����ω�[� jP�����ǥDK��Ӧ]�r1����tV�W��lf����\򯫋�����ӝ���@$��p:���p&��H�;���7(c�A�>����%,�̈́3���;!Ǩ	�-M�4�����ј�s�'���^C�Ji�2�Flj���&n�E�{�Z��ܑ\���-��.r�V+��D��y�b<@E-�@�1]&y#O���d��5���#�CԎ�� �kqv�o���ҤO���,D�<�@	y&�2�d4GK���` 7� �NC�S^��o���d��>�lDH��%�=�Μ\��MY̑#�"3��	��=�vF�`nS'G���2�r�K�	�lj�f|�Q������,7D���3��n1Y��ͅg�)�k�^���d�:ئ�F�%D�K/�p�ߧ@��A�7��hgs� [i�e ��m��N:�H�vd�d&�@O����9Ǖ��N�ыHFk&����[��6�2�Oe�|o�
	�O��d$��������e�&�_�{��x��w�7�Z�l�z�6
~��e��0�W,�0��S�Nj������eM�Z|��[��?k��]EùDMe!�ޯ�t��1�?6��
��Sa��Y/Dnm57��u'XճuH"Y��c��q�4.n��>K�:�mV��f#�G�}��vQ<�����g�f/e�V'rۿj�EJ ߈��ey~��ZX�n���چ�?$}��Bz_���R3��L��ĥ�����Ð�U,;��Cy˴�������n2)0�K̾պ2Oˊ1�K���A�("���=��ELk�%�C���o�Cʹ1�[����^S�NpoJ�~����:�W�B��H�>]���SM��H�U���}tӶ=��2'3��u'[%�u����C���zh�HFZg{���.�y���%��@�������Z���W���k��/B�l24��'��2G�y���7?��;8�:�nJ��p��Ul�p��s��*���p��$*ԫ��"�G�i��,�J ��M�25��s'���PTI>O�2(c�!��l-o��>�e�'ٷs���v�v��(�W3;/N[���Z�h��E2��ig��mN���dZ��Dp��t����m�p`�����I�U��Q�J��j��j>��dN�!�'Gg��� +�]��Gx�
�µ_ܨ�����Ա|D�r�*NJ��sg���?j�Ǭ�,9
������̉�ZmK:TG���v��a��`��}st��LG��,Vja�W�(������W˺��/�.�/�e�Yldc朳�3ifmҵ=�,`���xc2��Mz����`D����'_'������k�,�9�F�%��Ҕ�=�b�d�����A����#Dp��ܵ�Aޓ�4��g�j��KgԻ�
�{]��mu��@�.ҷ� �
WQ���Y�%�f���+C���/%+��*ޚ�m���YG������{�z�����?�_�)G|koW�jN�n��j�H�� dD4�:�r�i�R��"<Y����Yn�%C#�l�mS7�VlJ��X��`�8�g �����@�D֚Ms~-/�x�B�Aڿ��V�B��W������b9뎄�:��#����a�����<���o-S\?.-�c��.��7Gz �c���d�g���I �ㅬ�V:���!�qO�!9��+v<A|�k���R'<�U��pt�dP���#�O}����H��N^�LRlbb����;N�:��#�u�f���:i�^��gX�!h6Du��n
������Y-S�n��a������p'����.����[�F��Gj*��H�c9��7GY!���$�=˼�����"�d�k��y�J�O�o���&!��a��c(��>��9�Fdx�G�d�Z���s�� �U7l���_(I�Ir4*�cf+GP^�&o�]��d��(*l�_�p_\�a�dts��ݐ,�&
���ἅ��t[�CsM���n��ȪA̭ik}��kۣ?�J���Fvxu^����F}����)s���g�*��� Ї����P�1*�lqj��#
s�`�0�aX�%h ���*�<ͫ=��I�X��v �<�VY�S4���һ�ڕ�TcϮ�)8�G`F� t��K6������� �D�����y ��wxw �L��w�s�����.E��i�L0D���J�[����5��=�/c��5[�@R�f�מxp��K#A�Fz� 4V�醏 �/ש�g}�@KdG��cC��gqy��`���W��k>�{�����u�!�:�YًK99�au��xf��+�}���sN�B�� =���L�����S���A���^��Ճ���)��PE��ҟv�+LR>w�VM�?�v||ޛ��V�|lO�Q+���D��qQ��d}���*�0:	C=���m/�r�fn�.�:��tO���~9؎d6İ�F�� M-����6c,�^��o�V\U�i��c�:`ϭMt$m,26G���$$�,���(2c�a�<xHѹDZ�Κʥ]41��/�g���-���K.}Qڒ����w��t�e�F���#�&ѯ�s�$�K�����Qs�.�W�@��aZ�s�|�槕��a�ޑ{�<�0��Z�a���W!*)e��p�엹�@��酄�B#V�d�� �"64��nv�Y�S��0��Pb�ځ��x�8�ջb+��1wv%(��ɳ3o"�^�1�S6꧘�w�Oϳ�T��;�QȀoKeg"C��g�Z�C׭�v���697Kʱ�.}�v�H.!L�����4�o$���娌�����;h�\��E��!̅a����Q�;8�_q��­�	;�UbA�a�j�������o0ה��D���]�u���3^=h��n����Gq����+�*�ܩ=�T����_�����w�B�I	3?�V����[~��b�*4SC��6I)�ׇc��ao0\O� ���8�nB� Q� ����5�(�6:�z�<�J-$JȴQ~V6[״ܗr�T�C��q���[�׾}����J?���y0�$e�N$h���� QQ�3�-���jA<�d�M� �3��R������-%q�p'0���^������A0g���gy�j��h>q0����q�z��]�좔'�!R�p�����m@�AޢH[�<�ȭ�,�4q�C�E�Z�&�:��t�����eW'�/�_TԘ��-%Qה &�ɧ��+�?��������\ϼ����HĦ�9�B��݇��Y��9���=͖p��V��,�Ƿ#F`���>��L��5��S��,t:*���A8�@o
�CczDS�C�U�]F�?�"1�x�.��r�Xg=yY��c��J�`�8� ��̽���e cT"����g y ճ355p,m}�=Ǯ� ����{s���?N_J�Zt�{4� t�H��G�|���R}�l��ڷ�g��]}�-�{B���or:����uޤC�؆J��RXcr�B)�_�
�G��X�q���[����F�|�!C<�\�c�a=�1����-�Ò��o�*��aW����s� ����1Eغ<�t��.*���/��b[񥄪9�!���>H�B��o����~^C&��4�j8hG
T�m������ٹ:��$�*��t+ɰtݻ�b����7IҔ�*\�K���<Xٜe��_�xj�!�XEw	�����@�GЭS*U��"J��d�Ϡ}��w?K��v٨��˟e���+���l,�_ ��S��vz��QN��@MJ�&\���������~,:q�bk��R}�ij����.!�Fh�M�
�k��mƼ�'��|�Ѻm�W�UR��"�lH��r�+e��W��ֺjj��D+�^B!>'��
�*���� h����x(X���iO������{��|P�F0w�)0�ϓ$��>L4?�y p����8m�L섢@����n�2NJ�?�UI�l�3���A���C�!w���S�
+V��x�+����碒�+�����*��"��^��(���������*zt��åd�-/�m�)�}����<�g䜧��V|`E�<��,��� ���9uYЩ�B-�S��G^�%��kq�Kbb-!��d�5;�9��^~�㘘��j�RU"��[��q�.|_�i�_��g��M���{�6�t�=�؛Hb�i�:��g�����Ϝ�T�)�h���yx�ۊ�iXA/sX�Y�oU�Sl�d��[�n��U���ByJ��X���ޚ�L*S���Un�k8�+�rw�m92&��芙�c�z5w1 ��Y<�s��Df/Xu��z_ژ�(B0���Q{�rq	�����5G�Q� i|�U�L0���n�?�h|�Q襁26k�M�s�Q�w��6��>�ƨ��C��g�Qѓ�åǏ���^�b�
�(_�͠�S�Ӫ*��D�y�KX&U~�?|r ,�8k�;Sa��ٴJ��ැ�y�P�l�ق��)4�r,3��;�5<j�'����$_1�O��	���]��d )���<����8��8������*��N����6�ߨesPLY{F)$@�V�x.*�lB=6l"�����ۗ�`s+FK�kA��o�}��Σ��l'�kq˳��}��ɹMU8~��?@���H���+rw�s��,�N������cr�ִ\�C,��P�}_�����O� ��FW�o]�otC�����<bߙwtV�<���e�6`c�ncz��=I�o5�Wo�q�E/�x��O���Q�c�A^<���%���%2��krE;.�_ �Y�i`�uF>��H;�d�A��7b�R���U�=�8�_�9���P�|�Ie��'U��'f�m���b��A�1::��g����1�M�V�#dX���ЦB�o�^3���-��z�W%��ϻ�����a^ѯ8Pb@��ۀ4�w��)�\̏QoWK�Ko�TiS��cSZJ���W�U�A��"B�+!')��5�I�S�b���3���8.�6�1A�N��o�鋮W3��?� �����|xwwtG�A��c%bY��MXOXҞ�YE��.JM�[#�JA��z��@���^�g;b�6�Q�}w�u��ո�jLw,mE,��i����x���N�
H"��ר�?na�srg�b�!�Y�Rg�Z���;B Ӹ��{-f��dv�T1ʥ���*r�������5�l659b��[N9��RC�8��x��u��}i���cvu�V/�̋S�z�����q��Iה8SB��lVI� fi�91�+�bp�B���"\�o����4`wL��w�Y�#;5��Q��A+�,6�[�����P�ksW�x<%���92�	]�����\{g>�
���V��܅�6_Y�;��Mf/D�$+O�5��a�m�+�H�3���C���� O�6i�u7���R���-~]<�����	)�����"jZ���j���@A��c�t����f!�����~�"������M�VUk�$e�7ѩ�ig��s�
�<�S�G샦�E.�h��5��+�z�Ϯ=NL��2>�۽ �V���f�G��3R��1�Bp���@P)%�R��A0�ҥ��1�h,�G�5������@f ���^z���X=��RK_4t҂���=��y��O�h�P�X{"=e��h�xR�׋9'Cw�K���(�׽�v�Ȃ.���K9N3����kuJ�:���>!)��;�g~�07��ut�z�ԫ���=�ze%���r���r���RkJlk���ʪq�����y����Qe_1��]����h�gZ��m	-��f��P6��%
ΐ�G�X��=5����p�l������\)��eA^��l7�b#m�Z\{X���_�;JdF�y�=�5x�쳊�d\X�Y��ȴs���*ؽ���ß��r[��N̶;K��$���pGg�G����'�'Mѩ�e�:ҭ��*NR>Ul�噾0���ŵBَ�ĵ��~�����ϒQ�U��1R�NBj�&y�6Ƚ�*���и3*{��n`�dW�9yv�ª�p��ڳ��_2M(�F(T�SG�z�x�
w�P��wld�~O��nbJT�\FP��^S+%�l\��o|�rF"�#�Ѹ� 8�/K�==�B&�����(Ie��r���.�A?G���K}��e n'���)�2z���9&��Cm�P ��&��gS�pDMv4!��F���j�DE���ζW�^��ɬ%1 b��!<k�=O�q�N�]N&H���NDd�lM�[˨6d�K��a�6�iq����42��8j��q�`|��7���a�[r����ܕ��s+ɼt��d�"Ŧ� �!��{Ʒ��U���t����8呿0eb4��3�g���q�R)�ӻw-���Ճ��\��,�%J�|���E�e`'ͣp���|����I��n���*�+�[_P�ܖB�
7(��f|���,�Jh��������l��~�췢�27�֗]'�A4!¿M��R屭�Cß�d�^�T(�*�؁�f�kAۮ��'�֎�*���݈T�c�t��������t�d���93����x�u� SWFH�S�/������n*%�X���# �;y
l�.��6��RU����'�@�c\w+[��4 H��mq]��B�%917�F_ҫ�k�=T��D�N�M��s`E������&#��/�T-v���� ~r��{ӯ��F8��Ϗ.��{U���������7��-�W��aN�d "8E=p�
\�g�z�cTL�`r�Q"�q$�X1r�ry9�ڐv;M%_S�����S+9�I^6S2��2��6�v1X��mC�;��Yh �P'��gFLl��ػT���S0^D׌���p���zw�ao�ӽ�x������2��	
�xlO��)�F����_ô��s-��`�!KCPJ�	�{?��cK�㿉�x��K�@��e@fIs��/�9#���H�ٛ5�4(mH��?5@_�s�#'ޫSC�����&OQ)@"�$,L꫸UיD=b�&��Ny4"g�meY<_8�;�`K8_���������ɧulڋGG�7�8ҟJ�NQ�9~l{ڐ"/=������o��b�1��=/�>~�����Zz��WDW��:x�]'J
ר1�O�nԐGᜲ�q�.�%��k��U}�Z�_��2!Ӥ ��p�\
T���U�>���?�L��ۭ.[�����)�\��1ޟ������!�z��#��N��tQ���X�	�,Va�f�`�E7��������\���-؏���x��C����Ȗ��D~�ғ��f���2��|����q�3���U��=��?U�A���
�
��˱=�W"��]�@�2����vQ�h}`�( Y��D�ƪh|s|2�	S���Q��`u�J�H���Cb��z~�(l��	nLz	{,�i�2�i��8p��r ���z�̝V�T���V��mґ��QQ��6jX�=�'�M�BR��mm=�"vڪH�������q�jQ���� Z�Z
��.��FYB�>�+և�sIVc2�����_������F�J!��d�g��~�6�	�T�X�1��X�l<3����-2��%\o��j�r�o��z"�0e@�"
s���M(!\1��d� �0��iwH8E8Ǹ1>6���$�����}����n��b[�e��T��)���� �I5�Ѓf�2�9ѐ'��N�� �끢���lp�<�n��?�h[�aac��S���(�e���U<�X�8���l{�~0�_v�
e'C�':A.����)���z� *s��׎/mo��RS�6�G�Hj�`m.w;��Vnf�E� ��Q�SحdR��z�7���2�'���ۡ�d̛֟������^�{�ď����ì�s��g�M��o�:���V�g�g2}Y�h׮�j�� �:�:��%=�kyy�Ozg���,�a��'5�v/8O=�p<�L��=��n$�ڐ6Z�1�: �Gn��W�}�x��=_Jca��G>���\����Kn�'�w%�=��ԙ,&��{M^#AcG��8׷����<CjZ��V.Oa�ۚ��Ǯ���a���:��$�.}�*Op�́^a�l����� �J���+`-�WS]S7�����Ö6�D<�򜦑@9˥%Z/h-d`�b�-���*�UWj<��_Ku��\+�/�S���&�FM��5/�ž O���b+�aj[��&<s���`��ނХ&���痄9�!�!l��c���_SB��z���j"����vT�e$���o�[O7���< �6��X`j���[�l�p*�Ε��V��Zd�Ɯe�ry�Ź �v�z1���� ���;�t��<�j����>�+�����)7�W�3Med:@e��7�F�"��T#\i\z��M��C#f��r/�[V��tI`�>ru���aS�3sݔ�!e�z���#g�@RE��*�/PR��{´LArm�0�8�X՗p�@�߀��01���B=���%��ǭl�U��gGζ�2����lm��B��5��P��υ?r�з��tG���i���W<H�8Ugy��8H��O���G�Xq���
KrR(꥾�w�v]J�]\>��ďc��Kѓ�6�9�;��zM����V�`-V����ȗsc�&G��ڔ2���Vh�x��D��v�L�uY�%4�ֶ�����N&��-?�����E�wDb��&�����=�j�u��ox�IQU�6����<z~B%e��[Z��*A��k��[�A���i%�!�i��f+]Ґp�R�%�<�X�\`{�H>�$t@O������0��L;!���K������+�"�տv2�˕�(�Ac�,|�"��b2-�q�'',��!�X�w��WNE>��N�c�����Cѹ�o����s��%��S�8bˬ�V�A�12Ra��̿_R*� �!X2��� (9�=7\U�T���i�RJ�T9|��Y+Z����t�r����Zϔ�c$�-x�����n���-����oR��dp�9��;�[�H������tb�֪@��o���\[�,��B>y?�n��餗��(�@���²�$F���ݡ��x�S{����v;R�ԮNi����}匴�.�xj����D��?-2˩��}#�G���[2$\^q�mQL�`��k�c�ǧ��de W����gr������@����h��y�$�%�Fst���N���?�r�&�U���g��s<��S�䪶�<vO���
I'=���l�Q�r}��� �A�y���g���*r���#E�~��l�1�GVq��hk�T�ޢ�Ƃ=�˖���W=�p})�ȫuG8�0���ۏ|pJ��m}H�ʍ;ut*ن���T�qO�*r����7�$��8��>I���nO&��鏽:�-�}�^KX~�5�h�9���AP6���Q�3=�Q��Gl�'IĊ�5*UMvJ�8!��uw�����*�Fg��*��������T��)T~�`ָ��{�uA�p����ڂd�ҿh�����8T�^[��*+��~&	o��>��:�"K�g�;%@��h�!d�`~Y�m�oy�I�;������0��є��n�^/�z�Ѡ��4nrdl�4`��S��J�^����WtW:����&���b ג��#����w~�����O s��ưٷ�C���V�BS�*�9��٪����j�#����B�E0=�^�¦'[���+��I��Pw�k
�0��7����qDԎ��y�DNtI���*<��R����>�/6�i҈Th�>�n/_�%��
�$�/��a��F��t��h���W�vO�$�Fh��8��%���]��lX��E��O���VC�5a<dg
L8:���ž�ri
�؅f�����i�G0 ,��o�v��xO����/�(�>�_�W���;vt4Cn�T����j����J��@ Ȧb2:��!oШY�P����Fj�i�H��=�'�]#���Kk*R~;T㸛;3�S�M�����3�c������9����2�W��K��/t�z$!j�;������(�c���-.$���H{��:���&��M�ɫ�S+9@�h��e�����=O��p��d?
���S��
�Ğ��NA����@8É�N��@fҧ{y�+�FYÃӺ����8ۏG���
ډ�g$?���q���cL�e���9�L�G"���}q��k2u��@x�r2p���W)�?�y�pz�ָ���5h��͚7='��gT���d�fG�w-��qz%�~��#C��	������IK��.-f#8����:�KE ��O/�㌎H��1	ӱ�4֌%�lIY�3e�0���(���bT;��53S�_;��~��[I�W�
�ak��yGp�/�^����j)٠�:ұ��]�:Zx�_A*����,;�q_��������f��5�����Xح�T���0k`u����5�Z؋,b�_=Iic�־��ZY'O\	�'����=��di�iɕI�;d�Zݏj�lp_O���Jy���
���!��l�og���Q�+�����P�	D�Z@T���l��]B|#9��S��������v�����6��e�Q���?:��m)�%&�h�i:�,�9/�3�̀꬐��E���{K��p��[c�T4hAƢ1�W'���#s�"2ѩ$�=�Kq�X%��t�(��_�_C�p'?K�0R�O�@
��������x���9W��-L��5�}�����\[;�����r�ȕ�U�>����>z~-�Y�U���uHBwy7�������]`J�`x�M�t�/�}�鳯-cO���O9���g+��Q~MQ�?���5�2���C N��^�Ɂ��-L�%��o�n\�0N?e7Q��T�T#��&a�U����K��hr�>Ӽ��`�^9XC�(�ka���0��HR$Y�#����M�,v��Ǡ����K��ԛ|�:F�8�����nΙ��mn2#���nN�Zd��D����8�c���/��J����N;��~�N2�����F܊�U_	@
.1~�?���έ�N1��&�������t+Cn0�ls�՟�gWG l9!�7e��.������!����G�^��yB�.?���|���r�����I�-Ͱ�ga�H���)��f�W�*7��g�?�)�h�Y������nS\yqx�[l)s�`10Aw�Bv�R�b�\c�N<#�f�y'�M$�d��{<�:���$r�j����e��HR��J@<��w?��1�gmX"д7�����6g@x��e!1�4rm��'\��Q����ϼ���ԙ��1�hʮ�ҕ��<����v��0jv�v7�d��Z��;X��,��fި��X���#Q���vq�.#��>�}ZuʠJ�����s�Y}٘�k
��h�	޶|��*�D�� �8��]�.��m�}��we�k�o�s']
Q��0��#�y��8� Ms|wB:�(�"�eI:B���Q,LM
m�v��Ǜ�|Sj�J��r5�Kդ"�Z�R.|߷�I<TYS�S���S�kKpv5m�t��QV������;�aZ��U����ډ.�+!����J�H!�^P	N��"�]����s�%#_�I.�_�?(�F0Q��c$�I��},p@lG%I���cUdH�=�v}���R��[�����2[�<���[cw��?��m�L�c�Fo�����0���]�:۾��\��e�Lx�áC,���N�<���������G�Ś/
LA��=\I�ţ�y�KjV���i�����V�=��+9��e���y����C�����<�����y#��UbXԏ�I���S{���
���Zw/���4��>^�W{@����Ȗ��������>&��D��I�%^0�}�8;�o���`i�1�� ƈ�-�:;��+��V����ֹ��<5V�����E}�.*�Gv$����뗡c���<���o����i��5��X@��1��m0�_���� ʑ�A���8�����K�o#Y-k��8�Z#KPH0�1`:���C�:>N�U��$����>5��V*>�
'�;�E1��R�r\db���L����x����e�s����DpR"���	wm��N��>��6їм�@J7ь��5;s����Q��~�7�8�0�J�r�	΂�<4���i��=��5�&K�w+����E�M�S�^�B�%��پh�0j�;uq�g�df2��s�}�z�%�d���#ƀc��oF�:�w�U��;�)�-#��&��\�ޝ&��ӭ뺛��/�½������coJ���W1�u�������u��Eh����+�~����'�D��JgU�]�6��,E���#Q��X�@�β,]0t�@��6z!��������Gn4|��Kf,�V8�x�z�\c'��Խ�#�����xch����>��Y�l{bS7�#ɂ��i���{N����m���؎Fe�[�r�YF��'B�zwaV���E��ȥ������pV���>{������v��8�7m��'`��2/.���,Ђ�m9/?��'F�k�)#R�NFȐd6�W�/���L�h"�����M�գ����*�9�ÛJn�v�:�nE`*f3T	�.K�r˴3��h�H��#�KҟG)��z�'�D��K����Y��2U�%b�����$�'��R��<�(a�^��E����
�!�ߜ?����Q�Ŵ���2p̜��78����pc$Hͧ�~� �M��>Ճ%Wºx�(p5�	�щ�XU��{�a$Y`f�,�_�a�,�l+�t9�ͼ�w$-Z��и{h\>M��.Y�94�+Q�A}���pC�0�����cT5J�] pQш��4�ŗ褖��%��Jh �Pۮߣ'a��a���Lx�)I��z\f����9O���y��>q2�!�I�F��T��X&C��A�[��T	OᎮ��0���� ��J�� T��90�o�!p���%���ݴ
7����K�ݿ���y�w��i�@ ���y��Q"�<���ذ�����M�.Xx^<w��H>L�ປ�#�y�'���)��������ڸq�O��n}(�E��B&4p'�%h3�r;�P�;!�S��2#���x�Z��F��	����������Y?�J,nơ�Y��f �!�F_58��Yޣ����:5$
��М�)������:�\Z���:fѐ];~GOu!���"Y�܌B0v����ӰL�fn�c�K`^DZG�yD�.��vk�y�/s��tK�Ԥ�\S��ׁ�� ��i�[��;;���|S����t̟��h�7; ��l@��t�e�Ո��Qo�ѝ���M^�0�,2�ET�=��ɆVp�`���%�؄kt��o�s�(V?�zZ^b��q�?��=m��ƴ�zX����UMqn�H�.�0�v�qPnM��I�u~�K���OuPSl��pzq��Cح���_zO2���d�Y{/^��ɖ��yն�a	���J��E�QSL��д�r�^�8Q��(ah�"����5�ÿ���o�l�$@H���x��7��@~�ÌM��r�������,&�0{���Fy�@�x�Q��|$?�(��w�N�veo����*�%�,H���4���	_c���}�u"���
p�<O�Z��YὩ��T�̑p@E�B����%�˧�V�Xu��Y�u��}�T�J�D�o��+\��D�R���P��P���R˯�k�5���	����;z�/���	2�f4#���sNR��ϖS�3��� �����ڍ�^�Z�{{���@�v����F�+��#H�o�mqD$�Z-G7�'�mg~��m8�	�W�s�)���#��:,�Տ�3�1�K�/2�} {KD��	�u���]vg#�.%�7^��su)��Xp����Զ#�^C��u]���j�1)���D|���������O��ј�G�
�;3��#)$I��FJ���v. ���� Nk�!���k�1}c��@_F��Nh;Ȍ~�t�oci&>��w��㱜;�X�>�aJ���p_�"�=��ݫ��
��t�u�U�L�eᄆԇ���O�q��`x�
P{��!�ww�zUpkho�
!�ڣ�5�����~�=z�����_n/���c��v���Eu��4�6�*s�se�w�>��b����%���O�H�������8��ܞ�M�&,-
ȝ"�މ�O��gO��omB1^��/(M�[my@�.���i�J!<���±RA����ql����xf	9�C�����ځ�k�i�.��;f<4��:��RB�GH��z�Arg)���l���L���϶��l];�u�'���Mw���g$����v��J���I1zK�l��f=;g�Zd��Ť�ȇߛ%&��Y[M�d�ɜ��D,�ef�Ə�cq˪	8����p���D��E0�_b)��'�ؾv(lڣMj>vU�	6;�y�غ��縫�P�8N�#e������J�T� 0X��?\Y�g�8��w�1��u��_�dH��k�W�f�Zg^�x���n��l,p3�s~ЕU�*��]T���pA;�1ҿ>�U>��j�Lh���(5t�������a��٬XH��;��4E�nW�%�����hV��� w�.�Ao��^�TE͜�vi�JLԁ����,�LB ]ۙ�s*�6��U�U�h8Cr~A�L@��zJ��r�xЃ��+9~�=p������"����O&�J�B�%t�Ƙrn���*�s���d�5Yeݛix �CDV�������ސ3��b�U��n
���Ne��F59�m2a�H�o�����f>�Z�y�[�>�ȶ������Yv�7��v�D�Dp `�2{$6�ڵ�����BfYN���<S�BZ�|q�ƛ����^�)-�q �} G.٬.�^�؛�J�UM��Cb|�R6�b���?��i�����7
/�� B��&�4�1��Nu
���&Y�f���2���J�?q%�#V^����X9���d����sݨ�Җ���ֲM3UYII�"���-?���X5J���{��1^�>�tG�l �O���o1C����Va��;�%-S������{��bdUoڧ�w7Wjǟ=�r.���{Y�s�1|,��RJ�_���1�`]a�
�Z	� &�U���N3y)��Oό�ۺ0��[-�7�,L�9����/"�}bP�E�����S�t����b���̅��F� 9G=u��`��F;��1��A��KN	��C�9���,�*7B�)eRd�l?��ay^r�%X�ł�+��/��A�����#���bP���JE_�l�����;,G��'�gy)�k-e��XH��-�D��z�-8���E_�:���a�?1�[���'BGWC�WY��{c㢑�>���?���Km�$�}V��d��!bRfP�7�'5�^�����Pړ�M��Ʈ!�sX:�xV�Y}G=А��R1�`�IWm��RWLM����}�R��O��@�Iv�@:�V���V���7D���P.S�z�CNe"	�,�����^���k_^c���[���?�%������FnZ���^��s2�⊻Ք���f}L��,�|e]驎�m�l��$�|����n�+�O����3TNx�ߤ��;B�k�ȓRȑX��vM���k�s��G���܊�/�V�
����K�[�oEY+`��K�@�r�m�u'� <��aau=�����>���߀+��3'�e��U�k4���պ>��߯���ZU�T�P�g���I�U|4��p�Q,��b�|���;�9�W�z3��J�f?�|�S̼VP�E�p]���:x6_�6dO�:��a����^�	�^fp��S��j���Y/�ᦛBL�0�����#	4�> ��PSE�N�#�*�J���!��^�A�Xc���q��'H��7�8�)�'�m�
�Sg���ߧ�����Km�mu5ͷ���2ar:BZ�lY�.3���xt :��!y{ֈ\��˷�5{�c����˰�;�Z��x�Ɖ��_���&ށ+�`�:����o� /����?5{�P��pݵ���W��f�<�r � D)��q����g�)FH�����:�$Q��:9G��=�[��`�K+�d���'�C`$ ����g1$^$e�VwZ����fv	{�Յ%�n*��M�RP>~�mn��m���#nU�X���<1�]��`�
¹x��s30��D��"/���~Ј5Vc�)���	R�e悧���2�F��0���&6\#�| �QŖ)�����J{H�栜�˷�r"h�`o'l�vH���Be2T�ѻ�K�Ş��ݗȄ��%�69�g��6J����Ϝ6#���X֮�0U����c�S�"���!�@�2R�v�������Zq/��uz-Η՛l{%km��w��y�4BI#��<C*ne��#���aJps�.aЪ% �W(U"x��1�ψ�@X�����m��6��T��#�p�������s�oH�)#�Q&�����'���%˯������7�x
�ac}�jƣk�dN�;��p�eU�4�[^e�,s�^�����G L����rɢ�+C�E��a������ƚ��H�H ��4�MF^IW��#����K��-	�݉0��}��E������ ����1 /�6����ߵ'��̽Oӫ�`J����������::� �<����*�S~�"��Z�	�ļ�au��6�N�br�C�H܆Htn_a�z�B��8/v�Zo0p��4g�?�l���<b�(��S�
GMV����ԛ��Y�M��'se���W�(ݙr?���ڑpU]N�2
�+uZ#�oS��|�A���Z�%�-�F��W��#������iX���p1j;��-��4gٸ UF�a0Mր��9qٚf+N0-�y���[�� �=���\L9�T/�mW+1�V��l�&}��������Vʾ�+���<�bs;�v�QU��<�>�
h8�O�lq�9�)�Ѓ��!�w/��t�1��d�*P2�c��mQu�QE.�4���0���^�F���Qu�{�+�`��|��i �t����YS�{*0����=`U�$6E��j�?�E��x&�ݓ�wFJb,�mP5
���T ~/�����;�v>�:��z>�i-���q��2{����_�k�\�ܶ:�v����i+b?��L�q�[�uZU%g^�(� ȥ�_��W��AI�S�h�C��K�6Dܶ1��-Y]�����t�艬��2@%fff�����{�*�Oޢ�o�*ƣ�*r�}{�^���}[����$�KЖ)�������4��7��<d�$��?"s��K)8���S]�`��rʔ�\Y�[�����q4QU& �����Υ��5+/��}��;��D� �lu������҄�S	{��?�P���t7u����^m��pEh��U����9���?�5�b��I�Q"Mb���k���J+X"E��'��/WK�k@\|��]��]=N��/' A�=Ox��Y�+ FWR�Ak`��ݰ  &�2�G\ɹ���5\+6w��B=�\%�P��������(�\cc<�˅4R݂����t�~��A��9�f��s�2{�iv�cX�ƻ�,��,w� L�<�t�D�g_����VR�\�i\�1���5g;AG���:���h� ��)©�N��+�0zc���#�&�*j<$���������q����6�6T2�Lk�O+�K뛳� �^��#2m���7�9�y�8��z���C��E�3��'�\ic �X�u��2����t?����Q��
 ����	U��������W���\�1A���&Vj�u�Y�}�в���=��3%��M>��s`2m#�]������Q�
OX�l�{�|�����E�Z}uu~ز(l;�K�CF8�XRb�f@�jw��NqH�(C�>�m�Sr��b�b��ĥ+��-L���4����m�������iNr>Ǖ��d��o���_�S��u�����Ő,`��y!�1>RNܧ��劺G�)I��Ԅ�������[�m�5�i��PC)3ᙊ��S��(�p�E��?<V!q@��$�h%WJ����R�1*��^p�%k��ʣ�ޒ�+��-5��xb0u`��M�;�<?\��oՕ'p܎�.��4�+��ך�r�X��?3�ĲP2���(��zu��f�!�7�A�`/�Bn;��	������z��s�k��]�XCB7�δ`��07�-^�tD�Ǥ�܍%W�O��0F��@2"����F�_��-���*Ց���H���l�=�
���K"]s�w\zI��0]�HcΤF7h����T�'{c�p>�1��V�����=�<V���i���
�0ME���x��LE�v�t��p�V>�r�|}���^]��p�7��o'�37�[<Ei�d���I�I����6$]P^י�]���F� b��3�Y����wE񿾸LTd���/����ަH���g�����9��)躐�>��S$�]���Ԑq�Y����I�,�'�5Ƙ\k�����plQıc��m��L8[��p]���܋�Ҹ�s�X������~};: �cC�=V%z��r�_�:�	�+h���N�4ĺ��d��9r���ip���C�D�l�p�{���Х7�t��P�����x���?%V��e������JQ�&K�f<=�$�,�_�O&��|�9��&��|���\b	ɖ@��xbR0�$D�͟I��,ѶD�} �Ԁtď�M���C�,��Q�=�a���u�x�c��o�7d��j�S����5&�Q�#jBNj�L��Р�m?��R��l�Rv^P�6i���7_l�xgEֹh���(���\���U�&��̄�QS���cM���������\-]���G���xk����$5m8�3����jI�H�LN��d��2\��r����|�|%c�D%R��$+2�J���JOlV�8)ǚ��/A���~���9w\�q�qb+h�l@T�J��[[V��	*������.hz�k���KZ��|��Z�K}!%CH��9��~�sj*��l"���v�!T|7�c��[�qE�z�~W��g�ً��e��b
<�3���<�E�!w�����&�B�ː2<�X7��j�Qeo��wQ��$�o�-]R�-���ڵ&c �$F�D~�ɧ�����Ƕ����N�@J�E����U��+�M�XD^/᱁<G���k�>���#�<l���*����8P���Iq>n�ܖ���_���Gk��8g��c�{V��x\��t"��TO&��E �.VT�o"~g����m.��u�f�k�+¡4H=��i^��_�_h��o�6�<�����d*��o�s��ށ��=q���p�综�����F�K�B��= -4Z��6U>2�Z�������<�f֜�<J�#�
-��2fu�p�����7�ԆM��A���	h��Z@X�(%���0��ڵP��3)�3ަ�.��8al��J���?�u�tl[�ۨl�K�'Z񰠋L��wƶ@�~�eGO�`���3�}2[��q�'�2�SaD�D;Ul����^�oL�؀�l��FFT%2��SȆ$ek�S����3ʝ�S�hN��k�'�.�%��oW����zޞ��Q�X`O�W�;0"��I�ᶌdz�Xz[����ؤ��<�ۥ��`�ўT�i���}�e�l��H���/k�j�s�I��)\��2�o
e[�8Un��9�fK����L p�1��D�
�/����C&�(��q��"ɒ )R9����i۰��"��8"&��5�$Zs:��\��u �/G�*��k�c5��GÄ�����Ƕj��$��8���*M��,��X���]����*��I�T������ڱ��*3���!de����GV�a��C&� Vy�g=��M;���{�xTT��6��}eD�� x��+s�����p:�7���gZ��^D���B�E���z��h�/zڅBx�!�lnm-i�=o"�dׂ ���L�l��P;Y6O��i���L�{�_0B�8y�4o�?>�R��sV���q.C�8��ad�@��"�}rC�Y��OF�Р��'&h��w93�T�VT��l,	{��J3��[J#�W�|���NDI?3��"-�OΈ�a!<���V&?�aȌ`X�'�Y�>�}�v>����`ND����ae��
��Q�ϸ���%˄c$zK�aW��S! 4Z�y�H���'��JX��D�����Z�S�Z}�,��J�Kߗ]��5���#���f����� ��637��=�i������]'ݾ�:Z=vm���t�z�l�`x�e1��~�	l� �n�'���_�.�K0q�Y�le�A�8{s�BS\��W�+�k��R�l)����Y�߱G�WB�ǌP�#d���8{���	1�ks�lR��c���� ��9_��S>���}?$Z8&"�`������M&��n���ٱ ��mڳ��n��=ݎWSbA]��A)�	��pi�	w���������©ժs�
�)o�����KP䰀�}�^�La�>���]*6W|!6�B���d+�f��[?6�
a�P�HL�2��Å"�}���C;�n`����Y<�N��׵�~<ZS�d�RH�3��q�t�j,��	}��}�%�Ҕ(�3dz�7��|��� A�I����ޡʬ?"�_4��%4�*����~��y����[.8x�z6�P
6v2��Q�ި��<C����*�"��п�b����_�̐��q	��O��|������]��%m�b*��n�Ijo�ҡ�Z��i���t
\���n/�f�@%��+��
*�vS|i��ls�A�cB�K_k�k�ȓJ����q7�GP� ���b֖�pQ��RN�b���J�IN3=y�;wb�����Mk�xW��*4��#� Ie�Y@�xǼ�$}�P��p�j� V&l�=o�,�L=�`⟀��1��<Z�΄Ƶ�;X�c�:����)+��~o��V \CB�HU��M�f����f�G�́0:�`��<�s`��߄�q�<�����>�$T��l������땹�b�Q&<Ջ� ��HJ��QԄ���v�	��S3�>�(�e[�ա�ǺL�Q���V�0\z,�&߃��@��Z������&���8�K�3]� �Q䞊���C
'��ɖ�hҽ��$�$\����gl,Ъ'S�K-�	�މ\jՔ_f��B�64%gmǡ�r&�#�+L?�Ix���)�\��ڽ=�6Ү�@��k�eҾ;��t�;�a`	 �$q1<̲IlF��Y�6Tu�*IMǱ6�_V��ON�"m�3m9�5��s%�{d	|�5�������*�"]vp�k�kַIk��&U��o�)�a��6K}4��םD�iYK�+~
F�4�Ng���@%5;��u7q�+�l��c�aS]���ueB��t����+�v�Jn��ڨ���wYN�ņ���ot0�1O�/��=wt�m7�  ��ߗ�D����{����D�MS��1;�	���1#� ?�Y�1���S�."�J�YhN%(Q�=�Ӧ�DWUB��r٤Hh��t7�9�s$A8��`��n#�f����*�Ŏ݅�8�}gg���b�_E���tfVCP
*��j��"��N�y�tEG#{
,�?�("���hv��R���
'�7S�Y
N#!� r��-�ܻ/��
�F[~�Yis���+tin��|����+'�B���� �Y�܋!!�]۴`�.wS�<��͎s��_����o����V�1�4|%�y��7��d@ݭ��?���n����T����z0}�(
:�UXϺ�*[��������y��<��~7"��yo���Jbh� A��ALc0&�֏��Hk�����U�\��C=���2~8O%���P۴Qʚ���#5���)$K�J��ئ ;�a+˳���'w��H�PJ���A����/>kagNA@�˺���v��~f�����m���0`���>�h��C8q���A�0�"��<��VB�+"m��L/r��#��w{�T����V�#��U�1!A�K"@���-A�;0k�'��{I%Ak+*S
�e��� ���Y���W�
Gg�X�pYW�-MW�/ъ�f//�V�}���$k��g��/�6��;��W��;d��n�Dɒ�f�Zd#h�fu8�F�J�Jv*�c��L�	�
���&M��J��6 ɠV�g�WM��m/�5���k�oz �S�4�����!B��qt����D�u>��o�W�F� 1�!(١͝JG���ݟ�]����&�*��}0J��T��f.�be��� �C<������^�Ɇ�w��-X~�R`��%��H^W�:)r�x*X��T�ET��{� �z ���]Cw�4dw�Y������ܩj��#���i`�2�L�p���M� �1�H��v�_S߉#�.����=�O�q4������j(�ކ�X�`Í���HI�حw�Պ�;�`����E�±d|u�F�w^��-�-
ɔq��RxO�����o�Q���D��T���d���~���I*���k)�3��U���Q�x�?gν/�a�7�ҕ��q��������g�C���?}_ ��P������ca��;zEE���P/��͸�h���q��>�ݽ��dG󗞽[�>�?�Vwi��_�%L��B�F���	��N晾���8�|?�)ρ0ks&Ñ'ȫ��P �\�i�v7���ET��yȠ�0�W�� K
���'Nta?5З��S��PHv�6�0(��Z;G�*Zn��,Y����ͽ���i �B���f�5t��6�W�zN�i'��f�ԯ���&�A�aq�	r���$;�	ݨ�
�r*.z�w��_%D���@�{G+u{I��7.V����I�����=�9���WW������#d^?��P�9�"����zP>A�2��RB^�l��*M��fWB���2�9�]:��EO�t�S�k�E,v�����{ǈ�V�X27�������6�0Jo\�Υ��WqxS�b1���(��.xl�c�j�,��K�;UPV-4k���GQ��D9_��p4���@π�ġ��Y�Lc�&��oX.�S�4	Y$����^�	�����~� c8�M?*�mnz�Y)t���u/��k:���t�n���;�\�fҭOƾ`������u")a��>�j��߇��{���*��������������Mʀ>�I6/�
^�m�;P� ��Jy�Ι��%���T��è#n�o�6��]�C���K-�bN�ͅB�z4� 
�;e?ߒX<����� �r��G��,S0Ѵ�;r�SK�3���ѧ���S������Z6AJ�g$���H�������n���9|��:�H8u^qU�(�E�� {(�����C��o��8���5.��D�S�W'b6�#���G� Sd߽a��?�/@��
��%���<���]���ב�ݢ���	p\���b���L#�cX�띤+%�&nR��*]F�?���f�����t��F}����2Q��;G{$
N ��LC��ō�5�W/�(���U6U�?<�R�0X˟r�ݫ�=����Dϛ�;���$s�.�]�[��^7���P������Qu|�q�fqeTfM�\�d�N�l'�Ü]*P��F��ha~��!�)g�4���� �4Z�:�8T'�0ځ��8�rH�����S>f�MU�Ļ�{�o�gl�>#u-}Ɨ��D ��9��S�խ���"Mj�#��t�&e����1l�
��{�[��=W�10|�&����.�'LJ� �OL�P]�%;%�1��3�ίs�6�@Ы�)ʪ�����D���@��*�k
�5�1<����r�}EqrJ��M0C#����Ϝ���lHt�	]�Y"�qA�#����!;M���%\��K�]�jl�72�Dy5�;� ��B�֠�:q��
�!�&��>�B�),F��|��7o������D��e�~z���=�������A��)0��MS��k��mpC��V��)�w�(�4(��0)X+�7B
v���5Cv��Ŏ2����7�0�^�t0��q��2O�)���$S��<)j.�FqI��Q��^8Ik��#�x��4E�����ec�4V���j��{���2�7'1!oڠ!�^Q<r���\��QQ����K�e_�G�>`ظP5�?̰�[�f+�ǈ1{����_A�b#�b� ��b�._�W��s�S7_'����\hQt�`2<d�� 9@�yPQܴ��&�F$��	�vm�Y�1nY���),�C$�s����'(�"�����P)[\Ì����.���4��h�q�f8�\����!� �E�U6�h�q����ώ���e��Y���ܨ����Г�� x���XQ�<���>�mj[�5�%1e=�a�9M�n�!5����jrM��X�iHf�W�͍�Ǜra������*Ǻ:���ؾ��T�[c�q}H����l%�\!JM�Q�ߖ��v'�ɴg��߇�SV�A�vsJ���q�n��@E��lH��=���pԨ���m?i`�O������
��R�>��[��W�S5���9�9��-< ���3�l#�{���D��4��Ck����ٯi���h9]��+��
�����wZ~A�^��}��]U����A�ݣ�$��j�5B�i�Wֶ��- ���)�~6)i�8���z���=%������w�I&�	$���#D�Ax�@�t��oi"!װq�/T7�S�$�)'����H���6r���'�^�)�����!�%�<G����
������~�H|v��hw�u�j<텈0'{uM�oF<�]���iZLV�}٩V��a�t^�k�շ�����
�qKz�y3)i��V|�B��<Fs������������H�r5ȁ�����-��yaPMG����)V���|ל=T���S�>_�I1��t�\���ܬi`hŧ����� �MAb|�S�U8�҉�������gK��Ȩ ��6��7����ǥ��i�b���ݸ <|j(=�{ux�F��	ɥ�WɷU8`�slY#�;Krp쬁7�'�M�ȏ{NcX�)�6��t(��"	Q�+ɸ/m����+P��:~�r��ψ�ؙ(R(q@�Wl����z%�?�b��7�����l�J&$*fBs�$a��7��]U�sV�r�@;�{��J��
�˷$m\�tKA�([�:f��*C&�Ӏ�W�-�b�Ew�N͠����i���a������o������j`r�_BZ���#b�rϧ�����S`<��H��º<W�IN�`���$����[�Sf�(D����I�8ڇ�H>U��3޽g��u%� g�C�!�3��:!.�zFldQ<��Q��S�W����lL��8�����`d�w�ڙ�p` �@A���7��-{�����ʿ��w�[�%lAr;�9p�C��� <.s<�εF��e��>Rʵ"gְ:$���!����d����h��SIXK[L����j��a����<�k>����%��Ѡ5b�jF#�i��t6�lB��d�z�ҀMLdf��L�溳�e\Na&� С3���nU��v�-/:Y\T���&���6q���8�@\z����O�E<*R>Ϊ	-�8H'6��:��D$=ܳ�ᡂ� ���u��x���.��O�J:I)�Ǌ��F�J`�Ϻ��t���T�+U꒽�IK裡����`����`v�[CLd�c���>C<�X�Ct~v1r���Yu\ʱ@`�[�-��,c�!���IKTn
UCrV��K��N �Uu�yx��\�\:�d~��y���}���j �D�H;���3�J,��Q�# ���Qe7@�q�����ժ��篢�jO�V:��&��S��������V�����l��cZ	���QT��(=e�,��S��o�{n+C^7��9�k4�I���:kˎ���q݉�X�n�3DR��n��z�ow�r��S�����g�7bi5��������	]��.�4_���fMqva浢;w�����ax�
3�A`A>�5]���ء�?!��r~�]a]I���T�.��xD0�@~\���.��@l�&���y�1��ܰ��>��$Q�0���w���
Tpl��u++�F�� ��U�F=ƚ��Q�=%��B������)w�=Ac0\��EZ���Œh;�TV�U��.�d�;��:�ĺ|�,���Ş�E�aY���=�˘K��]��TM����#ڳ*� ࢴ)P����u��K`X�>/1v9P�I��	#ռҥ�+_i}������M.t7�9���ӓ�=�r~�2���n��K����>�V���z�H�0;{����Vc����.+hۿ���;\��^Z*�U�e�>;
t��YЈ*쳧S,);_Pc��F/;���"�N�:P��uEbkg�w�U�&ɞ� �������/������'���i>��;�D��V�O�C���f(,���M^�ɮ��fO��#�ݖl���nʘkvsN��"8�"��	��Z�´�m
�r�Mm����3Qx����9���s;�1P��"�K����� ��A:̘H�O�gr�n_�y�+��L�8�a0�1s-�l-��s��>&ǁ�Ax�����3��Hv�M�����@�.> ��B������uQ9B�*j����D-����m����W�Y��=L�Ք�����Q/��&��b�_��X��}{̟�T�_n��P}xZ�����H�T��[V�0�4b���a������m��5�.�ї������R:d�U�/��$��\>{��[�Q3Q�R���Bq1����e�wq��~�:Hī�R���W�(���|�E�u�:
	M�乾����n9U�kml06�4VΚ��Yp�5iCirI��YJv,�4�|��s�Z�x�m-�b� -U%7a�2����%=�����+5��ߑ��q1*#�3Y�$���|xB���),Z���8���ʂ�S��C����h�����Y1���V�1�! ^���Éŗ�l+'r�rJ�������b r���̢.|��tsG''�,��0��h;��k�U5�d���n��d�
��m2K��)��[��%��zB�?ǥ&��;d"���n�
� �����5O�>\[�\��O0�ꤚG���K���'aԁ
p��1�e�0ҜPhA��矜2�b��ֽ��12�ڊAV�W9R��c�/�%��G��m�Bf_���pu"���.W�m}�������qZդ��#EŽ��� �d�w����ǁ�(�Q=L � 0�U�����V�2i>+b��u}�%�0h��
V�:Z	n�<ozޞɯ2�+��/v�O�>#��.�3�T5�����A"y� r)���(!�k��љ�nWN�E�k����F�����s"׽ ������m��)%�G*���E3P�"���Z�;��qE�������5e���q{ہ�:c��gY1M+Fd�	�6��$�tP�L*�|8U��S,Ŕ3W��m3�1$��K��X�����bV|���1�.�G`��S���z+��]}���I���e�z�C�A�b*����RU�*�b�Q�	�đY�����e��/:z����*۽8���P���Db/m��6�f�����t0���9[ Z�b����cm��,��ǑW�xk�����'Rpkqk}��wLe�lFɗ��K��Ym�pl�x��]��W��<�Z�* ����<G�1A�|=I��v-�O\�Ut{�)y�J�3�2v0�w B" ���G�^,���-��޻tS��t�  vJ�G�5���:[�(�Հ���N�_����q�M��4؍��s��g��s��I�8+F���� x�c#�w��,��X�ݩ��j����;/�([�}�E�?��-u� �g2�B�v`�0qN7��m�
X��Lz&�N��o��,kjtex��J��[�X�r��0��>e3v���SC��!h�J���j����U��350'}��z����2���Sr��n��8<=W:��x��'�R���	]�؊��ݜ�B�<O�,5+���^���4as.�Gc.���(~��O�t��y!��Av�g��rc���7!Agv�;)�l�h;h6�qf+���
�\�]B�2U�{�7V|��*��Q?��)ʳ.9��!�r���H	�t���ܝ,uo���z_��5���+⟦q�Lj='��>������ � �_l���|�J�!#x���t�}���M�?-	,��� ���y����ӓD��7���=���#�l� ̒%���ݬ���e��	�>9=o(�ؠ�jeǒWL���0vſ�ցt���@����N���������=�84�OC�/��qO�����D�y6>Ȁ��:�ď�Aŏ�[�α��eR4� �7�Q��z)���G9EeJ�K��]z�rf�K��ٿت��Y>_`_/5�2�\ڝ�|l��z�J�F��}\��9�g��Ah})�e�rפ��c(������C��P,_�R&Me�@ f�?u��l>k�.V��/��C<�}����^D�` ,����h�[> �"�23�T��OG��)8-��}�����U���n6v�D��gJ�"����J��.�,h�²�$�v�� �n���QJ�\�p݈���f��&�h�� %�Vg��˾-'�s������ZU] �{ث1gI�'p@�1c�)jBca/�2���t�Q1ѓ���4�rm���X��
PY&�Ծ�__�;�p�VF��{aR�6=���i},~�A�H�'���U�z�R֞���Pg����#������=0�'/���R0Ry�v�K����`�#�����3-A�hO+��ܑ�\}甗
5c)TTy�� �4�n"��W������D��p�#Tx�����	��(	��yz��R���r���k��Ss���o$)-\"�SNZ��i2������k�ݤ�v�x���[�1�P^�������!�,î]K&�8h����.��Fg9�����#�Pƹ��\��1	�fH��+ߚ1 z���#˩����x�r8��gW�]
�cm�a�⢷�P�_��<Yz.���E���$S����"��5t2d�>��#��9�@;�}�sq��=�V%oZR�*y��W_��b��n:��Jؑ��R[�J+�^�`M�� 5�0�
w��~:=n;.�k�7D�,����E�i�*s`�%�PQ�n�=����P<�V(�h)^��ܚ����x�1Z;7���,�Q��C"��?���!?��r�T�iJ����rȆ�"}MC׼�RBFx_�ლ1荇�{2�+ pr������lWs������N3���o%==�ǗnB��<z��}��������!L-�Nh��pX�稄s4$4�J�y��J��F��,!9�����,�����=*��lgN��bf��g�3�is�cBoMS0s����yE)�AF7����+��Oyk���9LiU
����2ٲ����	���|�^.ت�����[A�jMK �6�.Z�@�?��E<!�j��a��M��FD�F3}]�$V��R�Si@X�L�R�)4���t"��Q�Jf�u����WV��8��u�Bs�PߘA�"�r���ܪ�C���Q�N��78VKtn�S̺�4r�co�
���y����
F)+��a.Qn�-+hH���[�aD	&J��W�V�Z��c=g�	V���u�LM1��ȗ �� �"9��(�2�v7w`�w��1�`jpF/k����x����ߡ��4S������Q���
�e�+������^�%��J#|$,��)ZP��g�@�cЛ��I�����Kw.HN\B�Xg�T#��BTVS�5��@�0���&V�B��_���<���(!}�R�,"X�~��+~�`	�&���;\T,�p_��1$���F�w��t��B�H�w����T��j�@p��U��~h�l}�|���Ƅ��qxI���q7�X�����B�D�է���[L釂(zKg��#t��/+|y=�����-VǇ��ɨ�]������!_�JOg�;Z�x�\��yh��\[�������a٥X�C�Dwl��Qe�~���Q�:�Y�Ð
�F�ǡ�se���������ŋ�����!#:� �d�>n�� �wbn���N��<����nLdK�Xm ���c��A;q�oǜGUh�>|֚��Ww���B�&}_d���$.�ߍ~��V����cg~����)�wr��[�dqW4��WY�f�`�S��;�^��3�w6�l��k�fQ��ӟ�����xZZ+X0��z7̭�B����!3MNIy�ڭ}}n���G��s����;ɵ�X�v.m;[YP�I��ycچ;ؔ��+}'���$�����w�ͼ�H�7�>:��;W꽗�-_��'��+¸�c��]�x���!�G��8��A�������_+��M��gx�Q��?��Ć��t�Arg�w�4ԍ�u�Wy5j0�	��ơ������o�b��	�i�XXZ��r�r�E�S�C.;��I����v�*�h����]r��N�fC�G�7�J����q�5V�e��SH%D0������2?Ӥο�����v�
����C6V�-����R�)G��fZ3(ڇZw���
5s��( ����d�K��H@N�S���2�X?�@�1��G#{y��Btü������Q6nJ6����*�[Tb����'��3q�������y��lZK�sċ *����<&Z+!0ӧ�a�RR�Zs٭2��b\�6����峤�8Xt���h��?/��9�ˊ�sבA���y�9P.�i],�
	f�5@a����I_U�
� ������8��6um0��N�]����h�u���	⁴���]��x���|-d@R��Bf�v�(��WG��%���;� ^�j���b��ҕ�����׺��=���c��^������˅_��i��D��R\���ub�R:#@PaCn��W�/�As�a�E�-���8���0m8����xe��/Љp�'���ς{e߽�m�����"UA�g/�R�f�R=��.����Wx�����<�MG�#�A��G��yj8m�g*�Z/��b�i3T%����*��"��X���}w������J�a�Ź��f�v�V��86�S��u ?���z����v��V�D�u��\W@�&7ܡ��xw&??B B�ՠ�k�PxL0����8� Q��B�W�O�iz�Ƽ����}����Xt�F�0�tm�_�pT�y����I�  ��������sEH�����X��f+�����G[8˦^����.�����P���8���f��O�Z�ym�������n�wg��v��Z�o]&�u"B��٤!>- )�x�������M$Pu�g��A�R�v����tݴ}09�}
n���p�/������Ћ����(�����m���,Va#g�*R��B,`�.=U�z�HL�HIt�<�q�z���gb6;��dV7�@=����x\#�{-��[q1��9;�N9����?��T?7�yi�=!��o�Қ��\S�h<�F�����N�o���%��MC�ˬ0;���lC.�5?�g0,t�%��0��"��"��?T�,��Q�e0�S#�K6�c6����+"o����\~F�@W�W�����s�(y���,�'���G=$V]��F" D=ܥ�}���,�1�t����!	*s�V�|��M������	&D�����U\��o�|"!wyoJz@#���[����z_�������Ԝ��)L�z�ݕ��'�p�n��7�jq�(�A�����2=��bk��u�By��C��_e�:~���A�/���m\E*��y6*w��B�{\�6���?^K��[�U?��]�xxُb!'�|�@���PMm�b"�����kTԦR�C�6ş׌�mA���ݭ�7�,VꙨ����΍�|M�R�e����)��.O�b���'�Gi��|8��b��U��w=KqK��Mc}�1���c���2̋J�¹鸢F��"/^VGJDܛ�q;OH��PL��@���F�� ����VmP�9 ���Vw�$�J�y������٫M톎]T�^S5�E�O�-��Dը#�I/�J5}&
z�$,x�Iu�9�Jo���Tm�W�vtC1�� �}��zX�n;8���[�ٳgS�V�緋����R�5V]�z�<��8��'l��0���X����ܻ���Y�u���c��>��W��Ż�E�jN�8��'T۠g~i����s.�'��I�0
= �/���-/(�Bm4J���3E�Im����'LO-�Н`@�_��ضrR���L�1�zXl���x�[���T�)��_�+���OU�R%v��B�CA��}���g���0#�١���Ͳ]C񷮙�,��W�쒽�X��h��
hD諀���C���1��5uB�%;qg�̉8Q�����Ⱦ�K%; -����?���a���Ɍ�4��(��$_g��.XX�v����8��R_'�Jޠ�?����n*KI~HV��TH:=jCζ��5��bc*���	��ͫ19��k�����a��CK��֓�x���&�Ĵ�[e�)�� ���SX���R����1�P"d�j�I�n.���йS���7�A�Q���4�4>�e;!��H�Q+��JYg6��V������M�>'g��8�+��y7	�rE֙b��I���V���:L<k{�1@}����woŇ��U]���^@4{��Y|���a��m��W����ؙ�2B#ـ�� ۨ�a�!��S&��i�X�HS�q&uDH^�ΠWlb�#c]��ct����δ8W�#�xYH�����[�6���o$�k�`�f�ʗ��xrs�Z9��M�v޾�5�C��:�G,���J~�(�.���x���a��x�5��;xJc��j�֑�ʛEI�nn��jz"ɼ�Z|��i�-��U�K�[iK/L��Ճ��A�������J��Om��$JM�����~Z4#�E���u��n�a�bKAl�T��2V�ox�o�E��s�^g��`1�Ư��֛�A�5�maP?uΌ!�Қ�	�Z5~m#�-&�,�ư�CD��Sҧ�mr�
CĪ-��g��"�v�[e?�%��!��䳀�4���74v�A)�DEE��*t�b�"�Ǖ�E�d�΀��2��� ���9Gb�J���B2�H�O�%H-C�5�ݵ�H]������I�8����D��^	 ��hc$�g�6B��]�|識U���+���$�� �Ʋ:@�,$���ܳh��O08 ��0Ï��x���8�Ń;pRD�������'؈Z	y?|7nd�w�<<����-�'����9�;S�42W��
��p�)�\^ƨ�D\n�ט>�"����?��|�?NU7k+�O�����,p��`��'S�Ҡ�/��T�U͠�T+��\M����
�+1.B{?�}��(��|��a"���﬽H�l�П~��3˛�.s�qƱ�R�-x O���Ye�a�Ssj�S�j�;���5�-�X��L#\�~��x(�>���}@<�qpɑp�UoM�/`C �M���RRaA!�sE����	jCB�6���@_��G=����f��i5���gl�,RT�+7��a�g�:VU�3��BӉ3�7������:���d�Ϥ�oJ�#���~Zx���7+���B�X�4�v�a�R��������O�)�Q�"�zP9�;��|�{��G��.((����P���5(�W���eI�k���8�nh�s�"B~����=i����,JBOH��s�� 8ei�����Zm�<P(H3,d��> ��������ij��#˄(�u�o1�$:p#��&WѼ˂�]����E����7 �E��*�CRA!�o���|�m뉸�R���������f �N]!oH,�j�|�.
�û#Vf$Rr���z�S7�� 3o�&�a�b�ء=Lup�N�6����i�f����[	���C�l�����ӧ��Q(��ӆփ�$�(?�Bg���s��Ǔ�O#�9~2��`9� #q_�.uL����a��j�ĳ����/���Gة7`��#��ddr�ң�G�*��H��H_}$����}�kb�҉B2��Yks��B'�?r>�I�N�Y�%�*S����<)6"T����5� pW��5ڹ &&΍���Z0�P��Bܛ�w��Z�_��� =1unU78**�
�7��`�0�M��N)8]���bDW����c��&# 5az�D����(��?w�࿴:�Z."��+�9�2���U.UT��&��~��j��3�#u��,	��3�H��[*��Cނ��TP ����E5��S�����2"��t1$dSC���$�_��Կ@�[���}AY�WQ���1�6�S*��oh5�c07 ����٣�F�y7�*���o0�0��O��j`�`<��=��e���r\���㤇d����r� ��KM!�$�fǦ�����W�B
0���Z���	uQ�U0!�6�eX�Y���(!�"�Y�45z��F��]kWy?�<9��%����E�G���:2��/`�w���(I��;��#�E=����(�c��L�AP! ,xr8����
�{N�1�?��<�S�W��kCd���&{��u��L�v;)?�T�+T���- �56I��ZŸ������-�0Z���K`� ��O��Kׄn[3�ť�,��Ѭ-w��=��\X�R�د!>Sr����r�k1�6lV�ut$����E�$�!���R�XG�
��f�C�𗨠?�q7���zַ5�3E�R�,`}ǓjY�npB�-�co�y|�3�r�4�S�A ��Nz=w��⃢��r���v���${��`���c��)ux��l^�I�=uL�n�O"�P�m�|YAnV�RM�^���F�w+4��%~R�������<�;@w~�� у��l4$��&I�n EA��d�-���ҽ:O�s�m�7_=.B�~��{��z��y�!\�ĸ4��u��}�W�c�?�MR%�*P��#����,���>"N4��Z�gآ �[���X�o���莏��Q>���j&V�\I�H�ƣ'�n>��qn�o�.p�Ƴ�I��3/��4��w���^�b�7q����M��U�S�g�'}��#u��P�:���>���ЍJ
6���<�<�F��%������l� P��.�ȇ�zeE�MY7�j�I*-B Lτ�
X���AѮ���@��u��~�L�Ub��!EI8�{�~�5�|d�(�Gh�y5^�^��]v|ƚ.�ْEƋ`�����׎nY"�t�Ӯ�á.8��(��̒��#��᪒հؐ(�/-R�L��Ԉ�ݷ��b~�9��\���ʂ1��]C'�/�q\Ώ3a�`����l��]s��}�����a��|<�U=�an]�����#��Yv�И4��~�����vL�j_T�/���j��������%g�6@�^�"�@��_^��青�"�HO�����za���C�π�b��,$�D��SNG����&�Ͻ�G��r��U�vJ�ܠ¢��2��C�����nU�Wժ���ZO}�����}�^ţgpU[� u���:��^(�uވ��m�PHQ���-���0c}�ŕ����������Nk��N��B�H�,Rp迩~��^>�i�K���xX�Zy|�,uh�WB�Z"�Cb�Vd{^.~�x����V/�4:ҥ�8��Τ��[�cM�sO�%eC����V��!@���#}�h�Ι8�k�Z4��佢��,P�P i�SȈ:� f@��Z`  l".��V"���M��sq�+�Lx[�r�����X�XҖ�+:sX�O�gX��������y`l}��P�##�Jf��3�Ǽ����;<���)��v��S�vSr��+�}���X����"Է�U�PG�J��!W��w)A"��$j��� �����[�*���l��Љ^O|A1�?z�=��+xQs�!f�Q��H	
�)|U.�v	�&b54,8Yr-n��Pw��� �ж��P�ƻ0�����:�K���i�N������ǰDa*��#��)Q������8��J��4����N8��m�p��1r�%^������R%�LX��_b����S̠}�tU8��L��9�8��Q˦Ө��T�Ѣ���q���s�{���Zyo��=�j͔Be� ����eP:2wr��:�v+9 ��4v�Z/���{�@d��{Z�ZqQ鱳�ϥI�6K�F!q�1ىs�f�Vݓ5LN�?:�w�<�����jS"������E�/Ob�ۻ͠�2jґ1N̟j�]5�W2��/��
�^�S�/�����9XN�@�i���Ԇ��=o���=}S}Ft �/%�u�xW_B#eR��g�_pi:���$_�b�����i�\�abwf�ܴ�}:�M]�IP<���WN/��E0S�nl� ���g~���g:�[��(��fa$��9����;�6 <�.�u�\x窱#@�tϵ@F�U@H��;�gx�_sJ�]b�(s#�v�_��ԼT4�Ӊ�a�P-~���G�8��ʨ�ƞ�<bmo���#�yo�{lH''��f��[6���&=Ht�*C��?��2�9�&;���ZҮ�K�q������h���6�B���U�q��f����C�A�/���h&�0��$���-s��PW��!(S�@��I�s�wN2t�*r�W�|l<6~�Nt�n��JT��y�x�Qd~O/$�a�#7t��M1��.����[>!bXxi�=�M�)ds������Ni��{	���wW �]��^XZ�p����2��>�����*%e���b���m�C����)b&��E^�^cfC�L����\���]���į4���E�&>�MBh{�o�ϓw���)��cy��"��q�7� \��Zp����0�V\�[L���Z���,�*�;�z�H�sy㬎zVX9}��L2�y�E��{-^�CG�~�T��'�$���V=ڟ3��µ�9�_z�䕷���.]��c�������p�tO�]�i��� H�Xa�������u�7g�`{��[����=z8r��4�ļ~��<��}�����������f�G���������'F���� zߊӏ)V��A#����B����7�_�/�L��@r�||�]�^�َ\��e�nm�k9�MC�D���qG-U>S¦��ځ�g	���;����L�{�,#�p�Z�¶1�z��Dg=���I@�}b� �ɩͽ���Q��;xmc�]2��%��3�?�����4�'��sw�f9�ن|��-�`�%�����.�g4L&�����pR:�2.�#U�̜��]BH�P�D'2��>��Y����%Zz�:�6��D��/|6���
,�o
CǸ���m�nbwpKM��>*O��mP�.7�w׫��UPWt���8P��ݙ�Fv����{�+���d�o��K�)�M�{b7T�-��ƹHjT��aߏS7�.����qYqu�B�n��9��W��UƋPX�;\j��-�G�A!�~��v�l�@��=a�e��c'*1�L�@��z�!��\�}u\j���7��W� ��%x�u����IhL.�{k��s��H��U���O���0�N��"��GK�;*���u~����GGh���+4���.���v"RgN�t�K3}���ޟ�@�S�*,#�uv?�X��&�L�Mφ��΁=����m��^mC�;g���C1�-�c���Ud�W�W�
��6�� �w�uq��V�j��E�^f�8Q��h�:���nK��{A��B.�1}!�U�1-{���{�c-�dX>C%���/w�I���d���k���?�;׏IO��yoЂ�\U�����'G�+�2�>�f����$žC�������0���&�wD�K���<�[�H�"����=��Dsv���版啋�+g--N�2�Lek!{#��������-�-�6���#�a"�"X֡��iX����/q
�eD6��mv��;R���^Ν��`�Q9�G����V�=̕�;�{+�"�K]7�����P��M䙫��2�V ��Oz㍝D]ޘT^�1W����QcG��d\����-$%_��&���a���X�.~) �C����B��p0����A#���>���4�GD��qzt����zc|Z3<�@�5&80���9s6E��zu�*~.>�[){\����k��~���8wx{�$��+:%��;t� YE���QE�O07B�	"@Xi(rvK����� D��5Ifw����K�{	R����G�\GN�}�Ɯ�:q��а��7q�xQ���p���7���$T��i��I��i4Ԗ��P��0�l��}bl�EN�P�fդ氂T�q��L}�K&��*�����(H�_~��82*�y+vK�jYNzY�{}v1���tt-����)Avh�c��g*�S�*:�`��KPvWf"�r[�}�4���������[�O��ŤWȼ�����ǌe�=s��l ?�v���xl�����S<3n�1�HA��{����ns����l?����L�7"����pk���� �j�rG��$=����u���m3SfnM#M7O{�*k�,d��=LGk�H,c~V��|�+���u����ɺ&��V��h�͕�$P���-�/8r�$۽i�o!��au�/zĴߐ.}Eou"M�(�����,��qK��P���i�F�d�B���Z~h�+����! ��Y�&�3��zT�A�8羐J�F஧��v��V�9S����ie�ӽ�m:�&��.��+� ��Nd�;��&��h:�@[�D�{�;p�~�s�����0���$�o�5Z
��Uy�\�.�j7΍�Ɨ�/�ԅ�M��y�]��Kv�+^4��<�d�QV�\<����j]���  �If���`��/#��(X�����n��N���2��+u��2������#|�x#��\�4�{�'V� �<s���ʩ�o�u)����=��ì,�Y����B ;��ʾ&��Y�r�?ߣ �{Ç�v-p���5*�M�)6��V�N�w(?&��r�Z���������N��A����<:?c y���F E����Z�a��f--pC�De�H�.��m�JX:c����.'*��?��n��Ps��.�]{}Ơ�Li�v�-��/��~�rB,p�_��&�$I�^/@&:���ͤ�Q�Kr�^�a�N�
j���W��?N��WN]O�Qod��?���*����f��K�a�|Or�9Ѽ�<����+�Q|�=q�hHr���s�I	�5�(i��t�e�+��z}?�zu!i?��`�IT��J!�b�A�}����@�ܨ�ʼ&A�- ��&�bhJ��t���qSm͛j���_q���$<uC>�LDވ*���H�_i����P'��n.��5[���k���V�-j
1��kĤ�yV�tnm;1H����EJ^X3�^��,���2b�o��V>|�
j�@�9��x�W=�;S�v�>_of�aFkp0����3uwD���w�����<.Xr}�i{K�c;��
�[u���e-�U̡IUx�.@tr͔��
���R���J <��GU"i�]��;o�+Cj$�R��U|��C[��������Gt%�{��gt[�UE�~���P��pcI2��n��d�K��To��YM�"biݻd[k�eݽ��i����t����h^]'e@�Q[��̋j�*:�)UOK?{FCɊ݋����jγi�xt��3C��01�%Y=�S�J�G��d�L�����5~��Ֆ��32g�qwz/��|�U�W$w�O�\( }���+���~$n.�`�Z�iY��VD���Hz�;����9��j]-�@i�@�,g����\ P�z&jo�yh8v�v��MVN��f���G�J��?&D���l��$L�	?�N)(�B��<�9�Qp��Vu��D`�8��Z�D�K�v���<�>�<�W �b������O�:х�N��v�U�B1hf�l��Ȱa�O�$�uC���`�,�Vhc�0;�0vd�+mC!�8	�:�ݰ�>@牖�S����%�;��R#
��G���;����y�Ul��E
�G�[�����ʀ�\Z�/@�Fp�a���&�Ű�g��Sn� ���I�ؕZ��i��5��Qk.����3v�)�Rs`يP�>ժ�8� ���G2�`���;�<���G{�η��.�,��g[:�}���}�Mča�E�%�ˬ�³��~��LN�i�5��b�"P� ����{ν1`�8�TYyU�3D�Q�E����A�3WȑB�u@���yfe�9�3i���_��}zt�F��Wn�YX��d�_m��pHzd�cˈ<�5�Z��}���A�;��6+&��}���+�c��T��J�M���	�`wB�D�ž���"�p��Ƅ��(ʹ�M�0��DK����A=�Xl�1�	�k��nXO1�6����v��T�N�,Q/��-�q���e���Ƿ�/�����^4 �͞�M�o-$d�����L��,�s�� �;� �X'��+5�Ҭ�C��pJ�M�p����y0L���(K.�S����^ba:����E�lc�Qr��)�j��qq���i���G* �(�~�D�rGL��/R���B|Y��;� 0i�!�=��3	���n��S�c��+u�,�����\�����v�� PMQ��U������$��ԝ��.�yGc�Y�����0r�p7��S;��ly�w��3��u)FGML�e�c�^��d��^��W�Ğ�ɉo����p�Ŀ|�`M����K��R.�GGj�FA{����j�2E��E#$�#�aC���(�j�J����,9���.�����h��ڟn���A�m�q��{-�H�uT4ɺw4v����k(�����ȑ��_���q��5=tp��qȖ����hs�Ͼ�=� `.����Q�L{Q/[�#�[3�\h�|���M�P�cz=J��?�����:�Y���u�%�Li}2�u��4�#���,�W��t�-��ʊ1x�V��\�Bg��|���K���q��Z�qY����\P���<�e��qSuN�Y�S�d�}+�A�]�U��u��Z���@��H�g4�g]ӱ ���Ģy�L`mX��4g&6��o��t��ˡ~��.묍�ZvG����h�ي���J���s��w �ȍuި��JYԶ,I�6���Q�HH�
-k.������>�sêXw},�Hh�k2T�8���I8��#��S��s3�����ե�E��@�ӡ/�ZmP�P^�wo`H��F�Go9Ԉ��dRv��Ns�9M�.+����VH���2��t�x;mĵ'͜��{�a��|���$[��
�q��[\̲־�$(���!�I�cXu�q����0���G���_�F��H,Qf.ҵA���7�V��j�l�#��C�;
�kϵf�d��Ó^Ɂ�>��	N��`�RÜu �Ƅ�B���:�B�nH�S�7[񁫆`�����z{h15�-��o{�bIu����,��t�&�)#�E=4�Vzrs�a:���x:8;ߏe�[�:ŏ㫺k�)|�0L�k�,;�M>&;�<nd��e�1I�$���Ud�/Uп�b����i� =��\>�C�"C�9��躯Z/� �h2]ڒ"�,B�q�<�96h+e��j+6;�QI���D��/�~��N��f�c�e&=�5`���G/S�1C[��L\y�K5Q�A�u���zv�(��hzb���8�FG����~��PP/2�����3�\Z�(P�?�t���AKT���ȀSz��k��o��v�U���%������c��z���#m�K�G�j�8 a:(�+?w��B���ɱ�7NĽoA�n���I��ٷc��~�:*�f��R�(�����O�%� RWD�P��`j�P
ݰ�TX�1\(D�wӖ���i��>#Ў�׷#>~,[��x��4�\�6<�?>�e�^k�ȷ��ܬQ�u0%̘�	d���.3�5��N��l|�ߨr��$�^��jgmxƵ�o� ��U��T~�D�*�hk�4\ҝ�!FeX�d6�f�^�liC-5^۲�wE*��>T������薤�YGR��F�EO
���]��Ckf��1���̔�~8������4Ҏz��tt��h�p��v ��[w�������Y;�Ǒ!�a� jE�s�Q>�Í�F�|v73�W�a�$,�;�����x>�d��)�])@bi�������9��J|�k!Z�m -EU���FM��H�3��<k���3�'�� �~�6q-+(3��DD�|�I�d������ܢ��)�*�h�Y�qBP��Zy�q0i\���U����)�ƹ\ѐ�G�O��,�A�!���*����Z,P��&~q����V#)�B����#i�*����}��|i�����iB^v���!�10k"��\b@�#���[�׍��B���2n�8O��cȲ�`�L�(���j�`�����E��'TG�������<�������&k9E�(����j���x�B�Z[n
t�f����f-+ekٷ�kk�x-`
|x�X+��ĥ�K�j�L��#�s��K7�����=����Q�^�x�%�DߩJy2ө��S������V����B�}c��5C ��-B^_�bkK�N�q��^�O��%�����]�|M�v>gZ��An��XT`�;,�A��m�*V�v��*�٦&���L
�]����X��� sSVO���4C}{{��!X@[rfQ��\y�0/��G�)���M�)�A�i--�=[�@�P-d!�4�G��`�j;�����nZ/E8�U9l�O�������`0U_�PaD�ul��:���!� �gL��[�A�Ī� ����t�[ �7������pj�Z>p(2����2m\"�)�Fo[�:�Q�93O٣�P7��y%�Ӡ��
O[�N��^�"i*\�iz�k�GfA%Z.�T�ߗ�*�/F��$P1|����T��&bM��'^^#���?�dB�D�P: ?�::뱝^N�Ig��̻Ia�ױ,�{,ch��d�P�.�QP�`�=Bq�1���G�,��A�̈́ ײ[u>��P ��r]��.4̯��_-�H�8z��j�>hz����R�c�poy�Q�`�L_.ʣ�?ɢ����%�il���������_��Vyxl�`MaT��2H��^	n:��L(�Gk	F��5�ի�:�T[7��yR�E|�z޶3p��[����ֽ?)�,R���H@�ʐ��/s�/N����$�\�����rw��e������X��P�q���5�Vh�6���HǄwLKZR����9O�ЉQۍ%3�F�Z¸�[������Qy]G���	�(���X�p"�щύ .�Z�)��a�O��dY`��%a�k�#����t��S��g���������+��MLx7�����M�8�߰�e�W����pT������˜7cȀ�:_����t�����e����z�BO���nhU���(D���Ĺ*����[�o�I�bXdo]t7��谧�pp�#� !��N�v�h����u�����v�e�!`��(�r[��A�se|�%�/�]�:��w:� �~$T�����橑 9v v���~M�J�6�����g���{���.�ҜT�C� �E4�)R�P6��FO[:v�����1�U ��{��0B,UuXco�7(��,=�WKV�^+a�����h,��7����8���Nz�"�?���n@K�AY����Qڰ2� ?�#��'�'���V�ЭiAx��Yf��̫�lS~���O��q��N3��L���>��4�����Rʇn�sDi�X���b*.[`U	rq�%T_�Q��|�4����w�R�!�yz�����\H0�vr��v� v�s!0q�(��264���;x��g���c\���J���*�:M�n����B��O��T�xv����7L���Q ��Z>�K�j�'����a���<�/>��c�i��ԡhh��#O�B^��5Z ;��)��g���j�0�\G���������t*c]Qg���!�T$�0������c��LLR���^���FV7lT��=�#.��g�˙H�y���l3Z�����taFh�$��E�ޥ�����<��nj;��9�5����v��������o�Ʌ���7���V����id,�(R�.�հ�l�	ox��t�3�}�h�U�&K�)a܋�W������f>��T� ����I`�]*�[�<F� "櫦C�Lx�����{5��D%�w�سN�+��*�0��8�P2���7_H �}6uq�mߥ�a{F4�ݞ��Ÿ��^&�`�1q��U�H(�E�@�b�U��Q�.
i��l'���WA���Ǿ��o4�O9EFqʐ�Ĭ4��
���r4��O+w�1�K"��Q����;�|<ױhb�@(|�ݎ�c�-�I�?&��+�
�Հo����f5�?���ƺ�(�%N��ȡE��鹞�q��U_�o_:��'�$�Mo�2��~�T�Kr}hx��#�:s��� e�=?��8�}5�0tZ	��\��I�y��:�?������Ҩ�e5�ɶ�7�d���
�<���ޙ�?E�q�A�>+:�w���n�4�8�ن�x1�M@�N��E�Yw���NqTCqu�	�)XD�91���sz�d���B�!�F����{b������b/-?���OETN�y�Y��I��-�@�&*�R#8����{�n�5@U=SS��}��6mE�'�U��\�=�1ѿ���)Q(!0JTU�!�[��8�In���6#�c�UAg+4s7�����B�tK/ۂ�s�wE�p��z�m�������M�2�p0h���״�*	(.�5p	9�OS&� �&@rH�>�qLD�6{u����`.IUI��5����	_�1n��T}z�i0{�h�z�O卝"��q�V�<�v
���m�.	$�r�(q�}���.��<�������	�xBׁ-5�LK��T�=DgU�+cݷ��'�߳���O�����!�Au�rNr��e��$��K�p��%D��w�A�j�k�� ��b*����q�*�N��T!�LZ�3�B�t����{�p����J�)E0�M=%}�Y�u��g�6��+tp&-��BN�Ǐ��9gNґ�[��޺]�xc�}���&UE�bvSE"D��\��LV&��]q��em~���v��"/��ɻ�Z h�eI|K*xU��^����E�y�k��e�~jb=w�xO�]m[:�-����O&Ö�����F$�[#j��c�'%mPlI�<�>��:|�{xšu+�q���)�A獖� Fj7--��)t<L�v-�V,+\��|mElt����3O����e/ ���82�`��� m�Z�R]�
	S���z?@,��WI��������N���[-�`��_0tl�Y��,����V������ĳ=C��)�!�5N�GTK.�_��N(B�S�g����Qh�V��E�>�2�hB�	�4��7�.>�KkE�=C�-~���E�"s��� m[x�i}�CYF��ݯ�B�_u^}U/@�2����n5�V�ua�$VA��O���:2�n��Ď�rb_���h��($��'4*s/'z�lHz�uI�AV�E�%)G@�#��7P���b3�8,����dC����bS�T:��������9/Q��ר�U�*w����t�8ٔw�~!�ҫ�_T��u�ȹ�$�P���6���8��6`�m���U��X�ϫxv�;<6�Y=k��qe�2AI_^����{Q�
��S��?vU���;3�/��AK�[Y�b�eMI1J��W�X����vUV�A��Rqh��9��^����%t�)�Ak�!�Q��k|���^�z�R�{�`��(�d�G��G�������6���"�0Te��1�S߅꾥�.$"ꋡ �����.��	(V��~�������<�WձJ���U�3�!�Zp5�Z�lqR��� ����^���{�l�u��,�v$ǨxB�,��p;�_����
ts�L�r��le:#��Lb�WI�M �!�K�k�-�S�Qs;G�^��&�-��ͺ/��L ������P�`�]E:��2G�� 残}��� u�C䩫�]h�hF�/�~+�ar�譻�)�G��Z���l浤_��RG��^O�t��Ndۛ���w���2��(i$.�u3���w�\=bz��Y�R-9:?;^ c���MUu��`�{�u�tN���sw*wO �HO
[hZң���)K�`p�D3��׏��7���I�0�;j������6����?s��A��Ot^c\~��#��8	�cV��G��と�%Ӣ��r+k��l!�9���'{J�;3N�}]*�ָ����
b�?!x���E��;S?!�����v���0Ws H:�k�����GIMA�X�����zv򿁹�\Wץ��I��*^��l�����w\y|�0+�#ʔ�$�#�#$N�xZ�'��-5zZr�����%�}B{�ǆ�Iƣ\	�㕽K1��ڹ]�:~����E�u8�N|���m`��d��������U:a��6�v��P:�~�����He(� �6�`1,�Eo��v��:��)G�����댳�����j3�d�z���O�6Ѳ*��Z_nWP܊8�bDj)���θ�
�zP�Η\��Am���ôE�Z�B���DI�[���$@ B�nP+���@������]ɨ$�o;�A���U���}!)��m� ���"fZt�V%����­����=UM�U���=�
�t:g���W��kT�D)���N�=P��d.i܏z�s��_O��𻅜p�IڗY�(�P�@��zÓ.�daku���:,b	�3#ܬ�׽%in����Z�1�Q����Xʢ�ߜ�v�_�/A�� &V��w��.���<-��C�������� 9�e�ą����bn��]l终�t���ׄ���Q C�5	\� I<��~�5�R������&��h�1325s_��',*1���x��� ���ה�Y�n�̯�6|����%p�؋�FP�2��X�_������  q������:�3�Y�ۗI-��m,?|�3M�/�l�m�+��)�Y/�}P����w^��tU�G!��I�*�����m%q#��n3���Rm1!�j8�!|�wq��ȸ���G�W���v��F"�)��q�"4�O�U�=��ݿ���%`rИ����0u����KF��g�@3Nɼ�)�2����5/�͢c�\����������?&��B,l1{�v��tzDɎ�,/��>�W�`y�3=0F��!�Ai�w����$��vZ���9`�[~�k}*���CXB$�1�`�'�Pk(�ҿ�N�4��䮖qr|�F��Y�[� �ϔ�%-AhGg{��
�;�Gp��H;�6�ǤDہ���B��E��(+#J\5�
��|�v]W9����	�O�*N�轔O����_����c3�6�Z+��J���m?w^�}�M��գ/�����i;۹�k�잶�q@��欦���3�u���t.*�0�%�V��W���s���<!M��q��L
��V�#��CT[XF�T��0���D�ԓ���Ց�~���K��~7����Յ�6_B�48��1X�^���+R�LI��ʏ�)�j��4�;W@��|����m��0�^��)e�lKӏ�T�$A���=��țF��f�^������.���$�!ϙ|'�*m�����1 
��'�zZ��C^��X[E��i��d��������I0�Q-0|�\RG�sY��!B��ĕ��=�fj,���֟���(Y�ϺͰ����)����? �4O4�^�4�O	ÔO����/z)-'�E��-">�k�z���n�wl'�	�f�o�;��akоe���s�c��q�:�~�	{mI�Q�r�-b�2�'4a����c��b�O��(\��g^�Z%�iPK*Pc��Kh9޲LH�����p{����bu#���_T"�63ñ&�����K��H@�?o�GLݍ�s:�_"�82ݿ(Ğc2��,vd�f5�_��`�\m�9��pva���ή����'���Bݯ��Ǘ�XxĴ�T
�\Nͻ3*ZZ��	SKN��B���6Nha����3��k\��ہ�3K
5Z �J����7�%DU�1��U�A��Rqú)Z���/�	�{��_+���y]��w�=<M���[�G8Hq���6ҝ;=��m�q5��W=�p��W"���p]v�v�뇒�A�8,�i_����Ý���aCK�+a,�1N�m�O4����jobJ�f��R��W�獠�W�|�����lzd�f�v�2�� !�~�?���mU��1�	��@�39�T y�<P{�r��A �0.X7m�7-��޳z�SZ�B=Z�ٚ"M�ѥܮ	�Vq*����>�{�1y��?���&�-ϋn6��b@�Y�"��q+��`��rE��Lx�CȂ��� ;��LvWF�2�^����3��Gk�I� �x��R��ѻG)b�eYB�D�0b�\�M����!g�e�1�ԅͪ j��~�~	\s�����}hJ�͙8~F�N�F_Q���`�����\}J����+�A	$�KlN���ߵ�PK�]d����<T/R�*���ӑHl�q��O�.����K�:�"��%}�`O�+��d��no�TGXOj�Q��gf�E�US���{ȥ^P;$A��/x=�e��2��E���a�<�8vL������P��{���?�6�i�.,]SŀVɬ��K��ZwU��d�7��8V^�̧$X��SP����d�]h�	d�*QitW�${��2��"O~�����3Q�oCh?���g��3��T�l֜h&�o_�A�7�%��w�R%��������R^�3��h�ֈK��m08�R�,�M��E�
�X��W�M�|�}�U	SS���!����/���3o�cB��u3YU�l����oǜb;.vE�,%��&o���V/��]skaށ$A^��o���G6��s�o鷌[إ7�-�j�̳(�Ƣ�R�Za"�ѧ�f+�*����jMM��@ZM���p;�;+��c�e8��@��t�
�"K��+>[l۵�;� �J�f:%��}P�0;��Dc9����~oM��|��_x?M������xw����*���)���Jу���x�j���/��h"�}s�͵5r����h�%���)�$�_�pIvE�nV#���r���(ܶ��Ǖ�����KtuU�]��7!
�N�8�MA�Ҝ�?���m��_<XgC���	6�E�y�}�iF�	Q��[�zS'4�Caǟ��8oZ��i����a�/��2���9���6"���?�e;N�uUai�Q+���L11|��P5gE�4T�χ���Vk��=�>�-g�?K�g��Y$4�:�9M�F c�o{n�쩮d ���2e��Zr�������^���1" ��ү����3V�V�]����.I��2�P������,�ex{���������j�-�W���ƴ�+jOʅJU*�1�|h��ɑ[����� ���n]!����2D��,���饍��L�ʕy��u��J��]��tzB�ܑ4�{�)W�g�T7�n\���P�i��K�t���/�I��y(}�i��H���XJgjj�qzE�D�lMF�س��.^)�y��="ޯ8
��*��a�/�N��o��0���+��=`��&4��&��@)KN5��Vvi&
1 ���������B��,-�GWZ���S p�pX7at�K��)M}o��~]'q"N��\ii���=����ﾜ����v�t���J2��@/9c�C7�������,�>TΌ��"��sJ7
ZM|B[��Ķ��t� IQG<D�����Q�b�s���>]��2z��R���SĶrK���iĽDF=T�ķ���.<��2��m߄#(����<��B��WTT�Jy$뭾f��]�T��'-�L�)%��JW����И���+��$���w���+��:��%E�>>�K�u|�i;�2x�:1f�< ��g�<��1J߱��a��,}�x#�-�g��Zxl4V��8Ӣ�w@rΗ_͙����g
��L!��՝��AF���ؕ��B��`ޔ_�ot�o�F���u�y�#��r���&���y��w2a �V�j�6��/gR�+~�?<:�ڹ���[�1�d�&���7�⛪��NU6���N����������A���x+q����|'4��ta�*��j|%w�޵^7j�%7������MH����םb���ZΪoO�~ѷ�/�l�WAc����������C����C:�x�jy��c�^QX+��$�7|-P�X5�|�V@���ée��|*���Ԅ�~I}�,�����b��y��Ua��rV���q�^D�s�zG��ZV������&�:�x� 9�Y,���\ʆ2�+Jᇕ",�ն��%ѩ�%��2�����Tk ^�x4>�[!��X�����d�-=��r��)(wI�W�no�v�"�����r��6�^2��j@߻�R�;�T0e�eC%_̤ ӏ/�d�#�����C�&�S�������%��FF����e�Zc�u�Au�R�3j�zqw��;��C�A{�V�7���2ۍ��!�,6̻��[�/�P�;��$i�cq�+p$��sx�a�[Q�����m~j��f�qԨ���ZA������^sE`x�"��T���-��geQ6D'. v�)\1�����hnz�^?�5RJ_��A���eH*�R�i�0��z�_U0�zj��}����A�-?@�?C��~�uF3�y���<1~_�o�S6I�^���� ���zc���mҘ���=�G�xh�zS,�R}H@�����Ah�tN��K�Gb(L�s��O�v4��Hܷu;�\C��9:Q��w��v+V�H����������
�,?�I$��?]<!�ρ��ć����c��dh���<��^�FI;żn:�D�.����Mb������s���X�ٸ���B6�[l�F������jA�yM�\g���{��{��ª27�uc/~xd�a^��Ĳ�;��!.�#/rG�����Ba��<�?� /}R�e�-��I��}���M��=���fi�5oB���-<�[��1W�lލ_W�vd��8-�<ǲ>���{�j]|��}N��g��%��91��c��I/������hۀ���h���Sr�;�r�{��_�X���d��5X�PF�,B��Q�J�3��9н�8�o�"9�e�a���ZV��S ��q%�5���54u����)5Z|2}�Md1N���=�S������|��������$���q<�i@��ft�w�9ţ���KZ�R졒C<��<�?���T�eT���~�ܓ��~�vl/���hgd����D�8�eKR���js���B�z~����#�as:���q�l���$��nB�t}����,gЌ��4.ۺ�]��ݖS����t4��ݥ�������%�^W��,=}r�c|u=у�
Pl5�������N�t�"
�)�{l=� j�#��V�Ƽd�[!D��L>��n�$i��y6��A<^��s���iH\,V1�����Xʠ���|;߿��.H��}p�c�,�g��O�$�u���l�`oktBl�}�aҏ��V&uۻ|�i��z�Hde5ѫ�d����u"�/Z���)�}������R��d��y�:��0#'@�xq?��5v�9v��D�n�̗��Q�#cp���eE����(�j�M�OP��//c�m�v�_�A+�~��{C �9�mW	�/�fa��
&oM6:smI:Sw�mW��6��*Æ.ѐ�Gl�
o��%�<��r��B��Ģ��o�h7�����|�z_t���
�^ʘ:Ӌ�:��O]��d2�<��|S4��Q���ܹ�>Cm;h(�J{d?<�b�k��
�?�5:#�Dqq3Ζ�N �2V��s���C� �垙iF����0%U���Ç�Ir"���j���,_e*~�E��ICF�k�Le�����AF��Ǒ-vY�� k��T�n�Q�3`I�N\}�ǒ�H��_��.Y
���wJ�*�k��f��L����ҿ��;t�ѡA� e�Tg��r�2D�
h?1��6�ށL5���'�/��zK���)Z���� ����%�Ն~�C!CY�������)6t�p75�� ~S�lS��}�q�ٰC�q����hnWE�P�ͪ&UA�{�$|��[=����O�{6�t��6�}�t�aJ%�6��$����*y>��V���Σǥ�ƌ�$Sukˠ�t-�@_�
)�df���H�S�{��F%v��q�~��T	�Ѭg���������TXV}� N��WY�% �S��x"�?�
����W%SM1�:�M��F<b2��S!~���,�������J�U~�
��%�3M@<gK{L6���M��:����+۸4n{ix��SI�Q#�x�eNO2?L{&)y���h�0Mm�^�E���|�H���z��Ȝ���.U�2A��l)���p��>���֑�!F_oZ���U���@޺n�c �[j`��uZV��YWr��C0ò��x�-m����
T��2ʲ��m�� 32�b�AWrÿ�	Y��4��E̓\���;4῭#H�{�g;i��F�y<8�£�"�tI�nEj[D6I �w��6��O�@w�T���a��KP6���
c�}��A�hD��Y]�ӮM�kF�F;�E\"�U�kn�(bo.��V�����½��F���W�u����I5�����x�F�q�G��Z�Y��� �k�T�
��J�P�N��X��P�W�U�f^�$����}�O'����W��V�$��{��:uJ|���.�S���������'c+���R��ײ�+�n������ ����W�иQ8�j�6�-�X;z�� �W����KqC��%���u�.@��%�lZj�F��n��8��D����R�4}O�%>��.�@�@����n�hSV>ܐ��!��*�;�EH�{�W��sAFT�SE��f_I-���o��@�ѭ�{*��#�+D2@�R>�A7+-�b��[Q����O�O���r+b��](�SJ�5j��p�%',��=$nx���Bj���xm���է�J���@RلC�ֳh�D�4b����J�jШ�m�(Mc��:��n��F�!/7R�1.rN;���~�[K?L��y��w!��]�)OFb����2�j@�%_���*�
hc���P����XaU���Ä����Vٲ��M�\]��^��tf�o�[���@�l�kj��\�iN^�
���ce�g�7i�&Rp���ur7����_�viX}df[�B�tg^@|�'c�|�;��Xv��(g�x�{��8
!gھp��d쀸�d����D�`�:��;🇬TW�p���D�_R��6���y�퉺��p_�e����"���{�[���
�������̤U_� �y��J�Q�e=�뺭��q�I�χ	�}y��K�@���ܠD}HU��m[�GMC��.�����<O�<���صY�S�q㏗��ƒI�9��<����+e�����Sү�Ia�
�!N��PO����賮��I ���J��1#��{g���mb� ��g�&��
 $��@��R�Y�L���XV-���@�4'e}�����ƞ�7�<�Ϧ��ܞ�`5x�8�姻n���^�5!FMv��B�+� H7H�%q�iԼ`g���������"Br5�F��B{wJ8��rL����CpAw %M/�Pm�ykˮ(2��Y�?f/��l�^5��.lE����.r�7��v��������	<$��1�nb(!�N ��3H"KG�uBʇ��F�_�+�oŚ�4�j�T��-	���g�Yd�qb����e}D������ɥ
��s}_1�\��i%i��u���*��(�0�!D?�f�D�B�J���Y�+��K�}�:D7�]�' ����Ӓo5֘��W�t@_���=�FF��i1R���<�u:�p7 ��+�Jd�ﭾ㎢��cg&N.k9�mƝ��y�Η|���~�����߃�B��E7���4 ��إ&�濆2��9�`#P�Qv����<r�9ւ�z����Ձ�����z�`��}9����I�P����H� {�ϙ�n��G���o�1�=��y�w!r���vx�-;T������	.jƹ�x�\Z��6˲��b�52����~�뤿��])�`qa�}?����~�JEa�֧���\~q���%��>H����
��Cl@�ͼ��1px�Km
F$��f�y�	ym�0)������k��JO�E�%gN����`��Ӧ� ���c�w�|Zd��htb�rt�p����f�f��4ʴ�Y���!@Z�Wm�R�S
i�\��AEx(-S" �[SA���m�
�%u��!�MY���4P��k�T9]��n�|�mҬ�@��(��[Z�ex}���Z��ڰｻ>��S�h��o����Evf�L��^�dV�*)��G�_� ;,�|�c8�F�sA̷����-n�D�sn���o;�U�q^��bx��0"������T�Y%�p�ҳ�85��I��F���a�d�/
,�R8'L[��W���=pIF��:�q�pI�wCi֣.�k����dD��~��/�?�*��D���<_IA�ڢZD��F�Cq�y07����A�S��tڇ8�d9��nDv���EH�C�A�Zk�XT6��F���y�?a("����`��V�0$5��$�$��V\��FCH9�2�"j�j��b��:Z��\Kzw�x�.A��aG��R�d}�l�Ż�<��ī�W�����q�E�띿���u��Vn:$�A�Bo�8�5�3DI��J�5Y��f�W��D#� �Ș���^�����/���>�?P�F�c��V)�:~gM�f�
<��X)z�O�,���)Av��1�
��z�N���m�-������*V,�S�������!�GL��u{<�u���m��"�\@�ȍDL�����xr��� �Y<�	$h2��=������B�U�q���0o����	8��? �M��ۿ��1~1�J�d&x+d��Y��]����h�.�3�2^L�����*�+�����\�O�6����j�0�L���P��g�{�������"�eܣ>�YD��k��!�A�[��7��T�qu+|Ys��r׸�J}Y�P���I\31ـ��0�ä��ۄ4J�o�nNG�?�GQ��Ѯ�3Ix���ɐ�).;S�ؐΟ(?S��ρ�?'�%os�n�=ご�<�_g�6��|�#P����� ũ�e`+SZ�޽!b;-�*����?;3M�u�Q��c��+�ɱ_Ĺ&V�JK�\d�xC=�S��q�/�n�A�s��gS��8BL��>jr��g�ѯ�w����'�w��z���)��P`O��A�Hߟb	�(u��M1���O�R0��+���b�Y���G܇u��m�r戬q�:�&����%&�� ��QC,�ZW��T3sdlM��˳� ��GS��4s>:-.�I	�<����R]?"h��oN8�� ��bSN�b\�/JO��R/�ҏq,!�i�`zH���߼åh4�� �ü*������as
,�j�C50q���?5��p�@ؚ�l.�������=3��D2�Ns��a�č���"��kt���D��G:ߍ���(� Y�x��DU�8�캷�(%�]�Wr�>�	:
:���U.���ܳ7�C3���=�&��&Cl)5d[s��?���b ր-[��f-����p�
�>�m.���t�8V�n;��xD�uQ���Am�'X�甩N=�#$�+@ULaN�4g�_�.��С#!u"����W-�[sg��.#q����\`X���c���؅�Z�b��ǣ͓0����<Vf��$���)���W͍՗�ʵ�eǻ�	��[P��U�s��J������ M�W�%�![�T#ǡ�*��G1�dG���5^��n�K�j�FD4F,��@)�%�^���6� ��Q\���e�Vb���+�:kٌ҅�9da(��4N��2)"�cK���=�K��{r��
f�h9>ߪp>�8���_�'�"�F�>T6�g�L8���T+��R�S4�^�P8bh|fa��+
�wy>)<#xF�Evs:-�ZR�Q_\��|��	ӏ�(vI{'5�m��x��w�K1�¼�0�G�1UE�_�����$Y�{�K
����˹Jc߈	e(�������0P�ܦ��C�L�M�;���(�z��;`�0Q�r�_R_��r�a Y�P���$t��-Ѳ��
�@u�Sf~`�������a�j��R�5�8��S��I�9;Äv�g|�ip�G������ܥ4��ܹ�(}��qf�oK��y����g*�O5}�z��|���@�b��V3�~�����8u!Y|KKW����&�R�'x�=D��u�oN�D�h-��]�߽<~N����,�&�j��󃖮�C��"w���?C�p��}�-����~S�
΁�U0=��l!W:�䱒"wY�'/��#��DIMڭ� ��w���I9��������^�i8? �S�sФO�p�Z*Q��KZ9�-�ϛ>���tL�r��R�-q�5[5�3������������Υ4�=?�� L��M�:n[ĵ�؀z=�]�����h�ۋG�4`-�P>��pv��ftDR��U!��=��n��'�D�v1Ui�_���lD�l=�9��;
7X�mƽ�cM��
c 7�/�����4[�>�1���Ӳ���1	�.P��1H#�M�0�mR#fjZ_����V?���:/�]����6 �Ę��e_:�������`�Q��ӛ3hB��5���l�Oł� ��l���R�v�	�$���������!��ָG��%ɼ����T*�$���;d��trg�ڋN@��Y�fq[�Y����;K�(�c�t�C��f�ű�b�ڵ���Jp"�dH����z�|ޥ<�g`�����B��:�'{�94_W`Dw�u�º�%�'��}��`���q��t��l����	��LF�̾4=y�֠f y�.��4!<��R'K��𞶷_���y�P>��&���94_���I`��N���{g���s�����m9�9xq�-�������,�9o�0e.U�K����r�)�
[��!iQ9�b��7���A �=qi��� ��CС�h�k%*�u%]�l���^�m��x�$����O*.��Clz"�"�%���~B�u�J�[r#�=0*'���__͕�A�m<�;�1/�$7D+����^Yd��,�g��
/�"yY4_i^C��?5&��Z�#W��Le�����)��d�>�D�-�?��w��>N�辴�Y8��HEl�TØ^�hm"e�-��R̭���?�!��R{��U�G�2�J4 IT�	�Bl<.Mc�l5����i(9�K(a�;���HP�a5�*!lɼz�Pu؛@w�&��!�:�� z2!�LK�� �P%3/��u��Ϛ�/g�}L# ��j�d�!���쉜At��QcjYɁ���4o�J���Q���V�g��sz�Y�	�G|�R��΄����ֺQ#�*cB�^G$�ώ���"����m���!*+���r0��8��������삭jD��m>Y��>i�������z%����)���vt���Ҷ��^$�m�'�w���R��9EΪ��X r� ���_gN�jG]$�x�5��Z^��F'��g��(;z6���b9L'���š�ke[䊨�YQ��N"2]Z6���G�@�ښ���v��B}���r���(�ʣ-�J%��H����Q����>��t��sʅmVC�l � Sv�N\�ru������^�zBo]��=c�<|p�EH�-�����P�:���oI���<m�0u�8��=��^�@�E��I�!�U{�p�Ѡt� E�u2XeL�RH�[T�-�L�+E�|��@
�s
1tN�o㖾x�d؟ɤ�:�gdw���q�z!%Nh8�&l�GG�x�QW���˧)�W�Nu�joP���τ�����2KEI��"�x܅���.�i��e܀��]zdkP����sͼ����r|�pA�/��I�Ɯ:Ҥ�U*'P��B���~	}?D��W!��LRQ
�����v?-^�뱍�:�a���]ө��2W�]0��A'+@�)�YW8�m��)W�"�	�%�%b��Cy�X����/+2�`�M��?���!����n���a�%YL�Li�\�#���'����Ma�����>ٌQ�؃s0��;�}d�$��<���ƫ��$�m�Am��
`�O�=�	�$�>
�uuȜ��:�<4�����K�P&��1�_�A+���4FD'2��|�M|W�?�7y�C{�I}c�=���J�ߦ���z��r�C!U�O��,5�������@I#�E�����r���kJ߆^J�o~���[�T�KD TQ�w���0Z@��l�,�=�1Ʉ�����OT6P��8;`���>QkŤ�~�3�t�FH�{F\�#�Gw�C&,d	�^�g@���ĥ;´�}���	��9 kH�>4<�S�0���sN|�>Zx�Cm������[�' P�p��ek�^��i�<X[2SȖd����YʝZhecե��8_Wϳ�˂%A�^��@�x�4o�i�;��x���1����%��C�+%�Y��{�ϛI�}Z߉��o��5������\A?)xm�`lT��Q~�_����mZ`^�0ˊ�]b�;�N��u����{�d9���"������]"�%K>���V~���"����
ibj��䨴�~�H�����)�M(�+ ��Q�e��A����u�Nɟ�-ړu�F���zDC�H�A!�4�*���f#f?*J�INA'���۝���W���Hi� ��{�O|�,��	�٬�w=�#�0C�[o\;���?a$](���~ڔ��e��,!�wklA�R��c9���mE,z@7n�С)�xy��9��U��qU��e�F�b��/$�3�rC�ؕT��L��9���"�a��m$56�`�W%�*E@|` ����h��#`R�5�K�A3Np���T+h7#��ʙ��:� �v��ew*{��x��C���
{K�b�B�c��T�R�$�w��`gg���C�}(���(9�
ƹ�� 8��"�@=1$$��u�Nyo�?����K0D�H��@���&���S�:� �.4� N�\���i<�-�W���`�]12l��j�{��J�T���K����E��vVa������.���.f�����ƒ*�`'&�dv}u�"��Y���c��(ΈB-��cX����b���@]:�,Ą��-�HsN�"�"���
�J�"g�Ad��~����n���lI�B+M��%��|G5��)y��͚ǃ��~;x�#���Z{ÞYk�N=�:���|�ɟ.,��,w ��v�`�B6x(�=�� ��I�:���l���;��co�5�"�Y��S�K����){�����5`�&k��<v�T1wgǙ�5��mw=y�\{���;yT�\H���]i�G�G�Ĳ�vn1�(��\q��.�(xf �Gb��9GB�AB ��;ǿ���{�`���0Q��g{'�1�X�o�]��feܒi���1э�M��9) +Q2����|����P"���F�ă�ŵN��{rKe�:S����dB\�60�4L�,ͤU�v��`�kd=V^z�Z3�x�X[��x�s�AmR���������l����M,fy�D�3�8i N��mGqb6STޅs���T����<�^�*o�ݞ#���Gu}����b�S�ց��(�7K��<�8B�ĥ�.d�(���K��������˗A�:�F����P�'�Y������z���%58%M~�2Z��X�����+;|��s����
?N,I��:�̒����IKH�-�*�B�h����g�E*��n���D>�[����������0.��Sр Xy������Y�� 9,Yf�D���
��亁�#���i N�UM`K�ـ�¼��5Q�ɠ�������7��~���%�I�թN ��J�^f%�
������.�]JR��R��>,!�S��Wi$P��[�oOl��gd�|)$B촤��^�*l����aۚt/J�34u�޽}�(���aR�?��d�ǩl���_6�<�b)7^M5�7�N�t��㵴X��`�u�O ��w�EX�����4�J��H�5��5��ɪ��	��k������W]#���DzȒ�P����N\བ��W����Et�*N�"Esc�����1�d�*��x��*PȪ ���!���E�r o�O� ~E~��L�.�Z��A4+ݻNM��������O������������4Hv ��>���z
�H�'=�r/�GF2���������A��fƊ�!�wV3��c�b�������+~J�k������s�ڐ�3�,6ʺ�(#���*~�W$�lI�hb��W� HG�g[e�zY��&JV�&�ޱ��eH7�>���[~(	=�#1_"�q|	��RR�C����t��k�m�,�S�Ʌ��qbH��s{*��A	jƁ����3�p��2~��1F�Ő���d�&ڮ{��U�d��m�x��V��D(ᗐ�C�C=�"��.��vn�Â�����B���
���\�B�����qt�Ʀ\D�f*e	.3�����`�}61�&V���p�ٓ�x	���=TF��,�Q!H�ʡ-|�o@��$��Y�a�&�2j����L�p 2s�e����F#S>��)�^$VT�����;���n�x�����$b���v��Ƭ��?*��y�� �P�p�e%<��k�7Z�~��T
8[�0�15
p���\2 ��U����v�R�O�aĠ<�z��]��dP�d��t�=�G<�5�� ��7�L5
Ju ��;9F�'u6�_�I�o��i~E�l��ԭ|�sҔ��l�H-�/�o�J�q$�jB� ?V_L�2�T�ʿC$=Չ�^,Tg���!P9�V�I�W��gV�m�G�~]ţ&�>e�_]�a�Ŷ�V�����������Zq���ӯ����/��u@?�<�x{!{R��(�|C"��	�w�f��LM��V�0��m���Y��X�/�O��ձ\�K_b&�^U"�l_��`Â*�,p����Nd�þ��a~�>??9�X����(;=��
8)IHT�$���w��|���H���G���'Yַ\�/V���C-����!���Q��K�!>�e��U�wH��J�%z�Q>(�(N$�9R���v5hzg ��z���Ξ6�?�&U�M�\�ڻ��wV!#�3���0��^8_he:V����]�}�ɉ8��{��ZT�JH��Tx�c�5~)�(��!�s�%p��(��!/�]��-�tq�4���j�7��6��T�ЧK�TU���+8<f�~������#��D3e8I�p�8��G��O�`,�Q%����h�Qf���g'f��uDnB��x��7ۆ����5
E���i�v��s��g����"ŉa�Lq�ގ�o6J��	Z�Q�o���݈���n߰��I�
G�fJ��"W�<贕�j>�J�BcL�`�Fۺ	��)�k�6�}Y�3Tb�����V�@��Pb��neYC�$u���	 ش�j�8Rb�}?�����*��!��LI-�Lh'#m�%�lB�L|a��Pͼ��]���5V�ݭf�8���.�j;�r�.�U;=K���Rms�������mJ�����b{��m4��4S���S�\xj��>#0$KNI]�>@I���І��H�i�|�P�^Qʺ���m��j2�{�Q�Jd�ᬃy�+�CK -6Riuf���<�eХ�&X�mt�4����p�6/��� ����ܼ�JdX������p�ך	���j��A'4X�Y�"�6�h��s����7"V7�s�<��ו܋Cu��qYd	�;������9�
�vҞ�N��N1Q ����c;
0�9���8� �� ���S���Z���ZQ��U��erv�Ǯe��M��m��=S�x,(����� � BU���R~�%�N���绨6�I_��
*u�?���P���ǔ��׍.�w�;]�O�z�M�Ӛ`jM����- of ��A�7W�b9"/�0Ap�f�w�2�Q��������Ħ��)���..�3����:P�q����l�eL��os� D��!�ϵ�H{�s�	�I��ns��S�Q�'PGoz��ƚ��>�7U���{Մ�+${`q��Y,�64r|���ט�Ǧp�#D�g�_Pڋ'�ƽ��_%Mu[I{�Gc�I 줿�M��v�[}}�7�fQ>_���dX����3������^���߮��6,E���G����j��6����dZ9��]9F��J�ms�p�	��"���$��`�23<��n���Ww���-L,I�3e����"ݿ��rE��Jox.�>�߱�u�p�_�W�J�A�R�\�g]o��eJ/u�Pj>/H��H�)�{l7�u�%P��'�&�+�녊;sω��VE:	೙���Ò����f�S
�B�v�e��u
�y�A����Y��[<N��pd��oF��7�z7��v ��q.�9���y�%�_	�ϻ�z��C)U�_��C�	���H�y�XFv��.�s��.���_o��!��N<"R)
E붴����B���{4�@4����H�\��K3lB|�{%�O�6򴟯m}<���X���ԃ�'��6��Ɍ���3�6wP�3j%cAQ�K
)_���䐿Y�$�I��LHcH���3��h��]r��|�v���69�r[��bb��1֊�1ov���[����Wɩ�h��[z,/4�"��U4��:7`���f0���WXϹ����vܺDҪ�{>��� #i��R|�k�2����S�4�}�,s6��&�r��2}���)A��N�_>���Ԗ�V"��o�{ڢ��R��̲�OSb������Aؘ�cn9yb���͚B#v� ��3c�3G]�mz�\be�|��=~n��sک���
��٫���py|(���dd��W@7WLb�I)nLc~>��]�o}
fF����f_b���vho��_��Y�U��;q&�sZ#�[	�*�CnX)o��?WZk���H��X6?/�3P�R͍q�y�I8di����D�K�J�<�3��+��?��HXo<_'%�9Y�7��RED��[��Ċ=�Cai�?A'��<�}I������Q��Ej98PDB�����y��T��of��Gͳ\vP,�˂oJC`h�!�(،���@���ղ��=�O�vY����,�ǰ�z�G�u�B5�b;����k-43W�j�Oyɐ�6)o=�Gc�z�E�3����!���C��b.�cAY��Af��|���̀��9ΠZ���!A�ԋ�;?�����P�l�/�j4<���\�_�0L-�'+����;a�6`� �mC����Ƃ m:��7=7;�X��V��ƗX�s	���,2m�M!�<�Ժ�6˓�<�;�]^�6R%�dދ$IMI��D�0D$�GTY_�	Ϛ��t�[���m|��m��' y[��O�p��ags��a{0IL�5_��Q�L������.S3Ӄ�~3���R�K,�Y��� հW9z����t�q��ܘCL�°��9�H���z���G޻��dc� бYq�T�u�#�]����&فv��^�]P����i�Y{�֩+,�u�0��%iF�+�`�I���!��nz��k}�Q�jZP��Dz����sP�L#�sS�	4����#ph�~��T˃*�b���%K�+�{��O�کL�k�##�{ml[b��;��ŝ���?��^L#�+=���O��1ΰtW�d	IX��_���/?�������طäf�E�7�\xW���(p����6���{������#a�T��ё�0���w��+�z���<�pu��\=�(!Hr�h�qA��W�TB��M��Iz })ῑ��Hj�Y	Ww�����g��p�ξ��8�-�K�D�|�@�@�@��^�����)�P��_xҴ�AJ�cP#�A�D��zF/{Gp'˳_�坬�/%BH�����db:Z썃h�~��療�	���D�]u�ш�����dU��F��M-�������U����D�m),	�ڡ2,�H�%e��� ���RҜ��WN�!�q��������fe�n=����M9�mچ:TD�iH[Z͛������%r�>z�x���-�Ѫ�ȹ͇���o	�=���1@p�$�Զ���7��ߐA�ڳ,?��z'���mo�R����&t
O������6���,��M�Ȗ�gN��ol�{�)�t�/�����ٔ��E�S���EORz8j�&�V)��t���IF[-E���(��wVB������כl�ͧO���`,��1tF���ǳ��aP$��CL*�
4H��}"�V��X�GΠ��g�m���P�lg��.��N6ے�xl*��Z&<��
XW�R^3#}]3:	��ۃT?��
'2�kV���kk��
/���-*�KY={�`K]gU>;�Pv��5~b좀n�`��2�is�W9V��X�䁦���vv(�gL�'/�NY<s|O���0��r��WFqO%��Hf���q�pO)����������q�Dxƀk#��[V���@�?���%�џ]b��
��ܑ��M�3[�P�#����j�h�@n\�?`w;6Y��_�h�D1���t!j:��?b�o[Oԓx��=�g0`CHT\�4�Z��������~�c��Z��\_�I!7|ю�����\@�Ơ^�c�>O��1=�^���zh�\�ep@��g_/ ���v�^�8N�j�Z`pV�K�n֢���̴���@��P5���N{���{�������,-�/q�(�'�����G~�r�?k6����QXQ?��l������A���^��r����j=GY��Uq4>���G����f.P�%�x�c~{l�Ⱦ��o�0���΁[B��
���r�(~�T�u�Į~�Z��&�HR�|7��
<I���C4 �xۖR�f��S+�1�_q�>]��U�Qw��W�ǵ):�7��7��83Z7�}����Կ��Ξg�}m,ծ�>�Ëu~Q�P��	F�p�Һd_~�D��+t4��~���wO�#�}rQ{�g+[Nٞ0��!�s��9Y�`���UН�v'$��^���kRO� �Ze�7B`KF($�U��@���7�����KA��Ga-VG��O�4���n;����#�U��H�<J���va���F�Xu�h3q�ʫ��$O��'e'C�sl�T�yD,�}e�{���~n,Y��\������� N?��{�B��u�J�Sta��T��B�)^d7J�<Ol�������ȩ7
.�f���ը��`@�$yQ�%�2��:�-�d���E/~���$��r,����la:���f$
�k�rq��]�]b�GW@q��<�Ȉ�~�R�#쭺+�%�nk���n���g`���,?2�)  ?���e2��&����~�5���d'��KN�C@k�=�Nic=%�A��i�$���%M~�H7�m�l��絽��K�g��bOAF�����If+ �"�ge�7��w:�|=Y�F��8�M*�-1��r#Ԁ�}!��*�y�9U��w�sl��e6��>���p�(^�g�2�i�e���6�*��;#�"p@���6���N�",��{�(1�WO�ݍ��#��7��
.3X�_6/�țn��*Sa��f�Su[��}t(���*��GM@���z5��}��w�M�h ����&S2")&r��U��S���%�������r�1:X{D�iEP�ﳘ�l���e^4���d�y>��WI��������pt~�x~BP�9@}��=��"n_�(���VGpj��܎z���f�%d&R�c�R�@��d@����1s�B��V�$�8p=1�����Y0c�\�]��e�1p�h+�GW��.M~m��}�/F��p�b�r"��D�W��O�o��5����t���^߽�f�Dg������� �Ca�V�k�|B�N�u�Y^��J�)�ysG����C�êK�C�h�ʡ/�r,&O| �^N]_��wX��2� o���5��jt䛑p���۲X`3TB��{��b��3��m�	 j�������m�`P���I}TY�B;��O��8��l�Ю�!H�}�}H��N!�m\�0�Q���nx䓚F@���Vu���3t�̈C9�ljoHȈ����l}Z=�,��n�B�S�s˂��:��F��;`���1�~�',��n��R��®ݧ��&�n�F��D��9&��� {�r� |�8��"��G��+�~'�Z�H���QLN4�%��nǤP�mOg��L�m�U�)���z̶b���'4mS��ʈ�w��#ދ��F:w4�$d�/�;'T�d�{C-z�ÆnR�=�.��`1�m�c4�߀����'x�r��*0�ؼ�tR�C����.~�@�H��?,C?m�uK��b����eG��\�^@T�;NfuD�۫��F��:�a����m��~-�d8'ջ��Dς�!sM�{�"�-���0�K>���Cn%T���� �E�} <k��{?��yN��Q4�9zdW]dGa�)�Е���wn{�d��Yޒ1I_]WcV���gV�� =��p�@S�1�T�3;�,����bL[�~ԕN@� ���'bQ���&+4S(;�b�ekΊ����ÿ|����_�E���Ɔ�V[YFM����~qU:����V���/�v�Μ���-l�(�{�~���y�h�I�Xl�\�9m�a�ĝo�.�|Mm��#�M/5&wG�
�P���jӃ�L���[�����PƜ��*�[�}&	�	n���;��?�R{	�b�4��¹�O�Ag�eO�:�e]V���M��E9�#>V�Sl���:bqw��ߍ~�asΧ3�'�u��L�_�6�x���]��^Cz��h$�gU:j��=GU%��OT���*kC|�� 5��r�G!}�}�Ey��}����=-�o��`�-�6�� �n H��?��9,((�膁���7�*�Ű`��I����'���^p�o��$v9��i
 �Rt�C�D}��o
Q����$��Ї��<� ��g#�B�ӏc�i�IG�~�T��eY�o��"5�����h�X\���4��:�d����1�+#�R�C����C��j��}���8Yd�'Q򘞍]�S|h�s-wb.)�QH��у˧�������L+��yO�X����t���-�sr�8�ha�Q��Q�qu'|���5xg�����?�Qm���u��e�1өl	\��)�t>��/ܥ|�V(oDI=�l�6��hVKw!!r-���P����S��E� b�9F�BAQ�+b �'U���9է�:�ґ��qI��1P����w�2�QS�2n�8�;X�����F�9ow
v7�o2v:~�t�D��$j�b��Kh�B2&�&O�$_`��EI���`����"�B���>8u����E*��<�m�����񣄫��! s)�k�C�K,��n[��#Q�d'�S�;���:n|`6�� )��e�G�>�e@
�6d�Z�Jzǋv���si����8m+L�¯?Q�����_<ќT[��T���i|y� l��b�
vQ$�H2CD����B����/wD�b�Pk�ĴM7�]X46%��C�bȟJ �Pq��ᱰDcCUs{X���"�]�C^�y��Ьg0����Ӏp�3vcqK�"�R���5�l�u�� �� �XL!y�E�}���9��6�����9 +J��b飜4aB��h�+�Q8�r�fć��ެ5(*�tRj��@���!�Ղ�������&vd�q1=|�XZӰ#�
Ɠ��4���aZ��ׇ�R��"�ک&�p��$!�F�Z��o<��3(����Q�]*Ӯ|X�GF��{3Ւ�mD����Ψ4c��g�y��o�6�ё��W\^k1�:��x�Gp|ث�����I�&F[d�n��Z��SIc �'8X�t�M+P9OE���li�d҂�����c"N��Ja�$I��� ��s�X}.����#�������1Mxa*��O�݆����s`�J6R�uU'�"qkV_k?��nF�j�X'R?>z�'T��]z:(���@�i>��Gf�&� ����5�
̀����wҳwj��q�sQ�K�C$Eo���s�P�^6@iy|�������TYM����d���^ˋ�m_��B��fz�U[�lY�h�X=Z>�}��
��4b19�n�"
�2�Q�6�X[���L�QMV����wD�Rw�6Vs��6���id%��5����^�֫�W��n�6�꺟O~�+Y���pE_3�����7u�̀�G��N���>sj��Fob"$%���3yP����k�#��m�-~	�H
�k�{�����Gmn��4�>_�v�:L��Rv�0Q�@Ӗ#���f�/��^�6���PT�4�"��Z�|9�]�'��$�"�}d<ݏb��)E����m�~b� !Hon!b�J�W�E��ZH����OԆ��m��;XrCa�Z�V-��Y
T���ppS �F��͈%&e��<	��*'��c-�=-��\*��H 
��
0��u���u*�ȍD��m�Lb��t��o�{��m
��2��uy�z
���6.l�14Z������~r�C
>�p��~���no����c2AOG����Q�+�̣&F�1��o?KpmU�tB�^A�1ĵ�Kl�\���>�S�Qfr�D{쬏�A_<�Jݑ�R�K!ѫIی��+?	}��s�@|
��#ŀ�� ��VA��"N+e6�j��Q�q(3�?h.��3k5e38V��J���.��Cj��9��m�8�\�Kkmmό�'�r�M\����wED:E4�?U�,cw{M�H<��=�I�I�L� �l���.�C��*�C�SG!�pa�����ڒ�`z�S޻)fT}BOg���Pm��DG�0���։��r�+�g0� ����B1�%��c��YC���i�,LjZh_� �#j��^Ѩ�+y�s��gP��k�7K��%!�ү3��&��K��jd�=`A�ƴ[岭)�����ן�a��C&��MQW*���� c���(�Z�ᄧ��i?���kX�nM�j6��K�4�2ҤDR�V��X�+r�p{(�s�8V����Q��o�v550�� �V�/�p��8y�_h2:
�
���L�o���|���u��3-���q1�Y,)3�����?@`Z��?fj���BɴBV­��S�A��*A��㤸� s���L=���Lp�ο)�7=wωgvI��o��UG[�b��;��t�m��J�����u���صg��5/"�A@�5�O�uS�=�+u�.Irȋ���>����f�>K��]��Q���6hx��'�1Q��`��F���~
fh��&�m��h�C�^���� �;��_U`�i�Ԙ}N��4 �Q�9�L�Qjִ�`VI�;pW�!.�F*6�J_�D���g�6���[u�(�:L�I��Ϫ/�+V�&�КK��a�`����ɽ3��g�&D���d&�0��ī6z]��{�)�+r�~�p��ג��8�Sx�y�$Z�H�;�N�Usm��KU��D
�1��uL�JOA|/� Ț>p�PZT�U���Bpԛ(��n�"ܺx�q�D���ǩ��RO_�n��L�n�|��mYNݮ4�v�S(�j�媄�H��@?�b���j9U��I�Y��n�@�_�V6�}V������g~��19|E��ۖZs��̃R����lPq�w������������iWѲ
��K��u���;T(+�{^@��#2�F����NW�>�� ye�c���fg�ZD�ʐ�m��|���
�V.��UKƪ�[l �y
�W5?��]0e�#��1���/1&���0�2UTK:n�̶ފ7*Ap�Dz��<1N�ٮ�B��^��M�rOe���#�o.�����Bj�鈵X�04}&b���z������n�ؙI���P��=�p��tf�$EFz��|e�-!�M��F �HՓر�ۅ%���B�����.T�P�ѭ-%��@6\�z?��/��R�� ���h�Y_Ew1ovH���ȴ:��|�\z��r��#�XM�"�GZ����D]sn������`E����cɯ#�[J�j��>��B��[�b�՘Ӕ�"��G�r�C��?cO�����T�����^�6�Q�3���*�AU�����s�΂�rEMJ_�O}�B]9kB�[`m	�(��������זYw)�f�6�ܔ�E&�D!9?wta/M�h_�6Y�M쩯�W^K��5}Z�R��7˲�����"��Yo�udt1΁�շ�dk��Ǡ�lb���r�
	(�-i��r�*�?٪@y�݁���r���,��<�0�m�؆�m�>�՗�<�D�zECD�ZP��K���dC�k@���F�w?���|������`bh�V�KC �-�a@������m�����a�#�f�=!�R�,!w�+�W��V��.�`R������P�Xu%4�}�i�f��L_AK�'fW��?:ˣ�;TG-60���~�X�1��_������N)'�(sQ�Ք5x���7v���~�"f�j<샹���U���O2��Z�w�_�����+p��'��I���$�]�j6���frJ�4&7��-&�����"�$Vn����Sę�y����k�\������!p���i�,�a� 7��g2|���rʟu��`����s*������цs�`ϗ_x�3�m���J����˶�(d��M �n�U'�y����˙�!Bñ��x-�͸��R+��C���m�T셗ٯ�N���JT����4)Ϗ�gX�8?w�+��Xc���8��I6ses���4F���w�D�Dd���LEma�����L��P�fDS-��RaĖr�a�q^̯��A̋��P�Q,��H���G):���3(?�Ѿ艳�"���qGZǤS�(>���?��2t�~�6t2�3z�GN�w�����"��p�,O�aŐ�BL�N��;#�r&4U]��f�yV�x����&��uK@�oV��J�h	q)T����7�@�bl�^�����8J������ꐴ[���������g� �ᏵOQ�=��q��FUc�yX��OԐ��=Y<��Y��a�07�(�����D�`7f��lvR|�g�͜�K����ŉ�i��I��`�I&�������Wg&��#��p��f!\�8�˾Sg�Ewʹ
�IlX�4�����kdf���V�V�r�`Pm y��ڧ�a(Ö
GpS,��s��j`"��I_TŪ¤X��	q�A���Tҁ��B5�r��?Ķꘗ�[u��:�t�P���{g_J}�\�X�{���dkT5�`$vv3�'�UT���N��Wa��M�띶��)0O}O����i9��t�T�g�l�U�*'�.Gr��3}V�g�|Qn6�ؘ(_���+��� 7V SDJ�*!r�HU��t�W\�F�G��2>z:��Ȭ�z
��9��o��]��tc?�7,��*�F�e��?����3�����~�R�M*�e9h@'F�PՑ���1�{la4��݀t9s+��`�Y�j�f�[�A�k��g�n,��
��`��1׍�-j��-	/���2�G2#߫Q�4	\.A�/��n�vS�zHm8�E*�?W;�pǽ۽w��5�ˆ�rv�PƷ9���<9?�BMP�g���c�HI�>:��^IG���G�"<${����#�=X�T��>)I�w[�B�Z�#]�������p�;�zL�-*ډQ�׃fB�9��7��kb-��2ףS�x"8�e�fvW�a�_dp<�t�@l������H-��<�4�6G��������ڷ�y���DݯZ��Ae�+�9�ցC ��fSɑ��3@�\�.L�V�n�@����vDc��텝�G��/�~҆UD'6�*N,�)�҇ ��U�������HY���b��[����"|�O,���]Ɣ4����wu���*����ŃE�xo���'��##��WĢ��ya7,=�X[(�����ui�`��ʆՙN��Tl�?]��d�Z��b<*� ���g`��i��](e����j��MP�$U*��=���Nj[�Z7�.�<��Q6�F뀆�ᢚ��������}��y��X^�n��z��P�/�[�����m7K�Wp:�� �������ꤱ8��`=bE��� ��ΐ%3KNV��� \,ށC�_µ��t3}�S�X�,d3�Hb������UmМ�*�X�V #��q�E_����X�oL�_�F��l�`�=��;�0W�|țpcD�AIj�ku`���x�Ӏ1��v�(�\��?:��D�W6��q��*�9�����e������t�86�Wab/��(��g���So��+�QT�G�KB*dga��ŋ���%T�X�UOo�.�)�#Џ`.W ��?!�M68�(~�t��ռH��«^�OCˏ���m؞��� z��F'^j�5@ll(��+:&>�-5��yX 35e�@��9Z�~�X�aH���D�?���N=��!2�����Y͋\d�V,r���� *={�H�*��ז�[��b�E���?�m��@#9��D�ջ�y!5i�ogr�r�K����.�2�+��fq2���蒙&6itΞ	t-�tș��x����C�W�QD��u~;w�aH��i�mV�� YY�)YUћ����;l瓠�@/�0�w��!/�(A[��we*��S���e��/��쎝Sp�C��BA�g�9F���j���t����-=�*�ʕ�$A��gI\߇	U�t��ν�K���������
��� j'�nx򳄑@��c� �##�;�"�qLY��Э��eF�쨡��`m ���P�B�Wd�Qo��zVz3��k<�rB?{PJ�p�����	B����?�)uK�`�Jˈ�p�N s�Z���?!l��	t��梭�R`��������2���i��U����E�K#&��1,��z��$匬ԓ����v9�ã:'�W��X>�uD��wdY>�^���"p_��r�t~����5�[	-ߩ���|i�Ln� �ycs�E|����V*�`���h_�6R1,uZ�C��1�2D�"q�G���~��qu��kڋ�>�B�ka��u�S���6��ω��Az0»����{�/2'a��vmP{���|�u�	zF�3���P���:u\�%whv)>����2:����HC�?Kռ�a�T,��AG�����	>$`/��6����勨��MG�KH�J���
d���~�l�'_i�'���mR�F��ۢ�5kc��`�8ی��o3ߥvీI��fR7D��q��3���ґ��Q������ukյ��c=����nƻ���i�B�������zb�>�m���(�U�(�#����<]0sդ*�G{�]8	I���}w{�w��${mف �o����
鿼[R�G��4&0a��\#1PH��>����㹓C<d���n�E=���	M�ɮ��\�_�g���f�)߶pH�޼��қ>\���ZB��Մ+��fy�e��|���I���X��{�ÆŊ�j�S�HPϘ��d`�����f�lm�i���Y3ՐAx ��&��S �>��k�0[�	�3�^��ӱ�D7PA���j�҄t���9p%5�Qd�Ǟj��R7���d1���G-Ôc��"��S��q�#O����MKkq��m��:���N�G��~���J���>ۈ��+)V�kJj�B5��ŅP0�[rQŕ���W�h���F1L.�8���,�QJl��v���B�#U��:h��<�f;q��YiO"X0�7��'�h�|���xE����Ve7�h�����f6�n������k�oXZIb��OQ��\��������##�����~o�M�2�7�m9.�9vT*�1`��4��?p�5����^.'� uklr|@���%�\(w�GFL�<iӏ!�q=�nDŉkMQ+�9P{,O=g�n�S"��y�|e��m�Mb> �=S����y���!�V�(:>fy���E��5��)�.D2����rV��n�s*a(���jB?��H�Ð�G��j�u����� !���(��7�?��w��c��̖�^�W�Q/���;7md�|��> 1gZ���Z�c�� ӧ�hwL�l�NF��\��w�w�ӢY��y���f,,(f
��� ?����rxiS����C0��ZI���r���!:+�6�j�4���Q�P�������n"'��f��ɍ�l���&9�ڤM�� ����_{~મ��K�B�P�㳚������D�S�J�uj@i0:6���1��Z]�����>7��\��\�&ߚ��	������*�p� ��W�Ba�U+RP�S5Կ�_�A#]��WR,@}��:0WL����Ը��.��%�dˡ�$Rl&^�v���Y��
��bdicG�~!,��i)��&HA�p�~i`�"�+~�_Q�!GZZ!���DV�A7� �b��>���#���Z�����������Ӷ�L�kiuX�<���ލ�`�����fnV�f8������u���}Ԁxc����{0�629\,�;�|hZ���yi�K깶B����k	UGl�4cY�S��R�2����K>�5)�AC�������p��K���ǎ�:��ģ�:���DdL|��`�C&��/ ݞx��D"i�.?s�|�ZY��8<��%��#u�����oV;�g@0y|�dBR4��N�_}�q)񁂒ُ�řϪ?�D��;{J���Z��<���}6������`Wvw�;�����5ԗnR����7^�A��"X����T.!U�(b�t/���F��TqWJ�9A���(r�������]��^�t���<Q0�����"�9���H��r�Lͽ5�yq�~$��+��
r+��}L��8�H�l�.�yP��o���0mߘ̴��$�b "��!0�?���J-!,�5޸H��t�-��'辉uB�J�C^�9���a|��Q:qD�JY�;���1B���F��2P�G5&�- ?L��r'L����= ��ֆ�aJ��o}���cX���'��';�8�̆eS<����u��a��K|@ڼIX�z*C�AXɋ�H���\��m�̆Br��cA�65?�n>8�	ߞζ��-�e�v���9r?S���n?�Y��L@�{���ֵ*d�Im����Ǹ�8��׬Y0rCl{9�/������0���׭���\��O����0���(cw�eS���O<�p�4��Q��ߐϲ޽�	H��ۍ��2ߐO���B�\+���|�R2�|,k�J���d]�ļ:��Mcsk���G�Q�A�Bm�����=�)�$��M3�=�0�>]6��y����t4}2B���A##ä́��]�5L<W�f�ϿW���Q`�K�s�:�|� ĳ�8��W%�t�w[WYIK-߮�����L�L9������a%] F.[�,�Aƶ*8�1\�(gvou�C+.�:e`�~�Эc�<��~���A�TE��)��ȡg�	
�Y�R�:E�{�UZ�_��oΎ��`�<9Q���ހ"|�;�`I��*;e�	mcG#ۛ��l��zVl�HմR˴Hx�֥�4ǯ=m��J����|"�čƒ$����*����/l����dv�i��X?�SGhK�^T.fe�U��uX����n�53oE��JO�G`�� zu%�w�[Ț���E�<Ń̫MaR�*-�ΧC�}� ��әy��iL����|+$�����{�g{L��*��i�w�`�"��?���x�:ͤȀ������	Z���3�gn�"h�Z^���}�����a�/	j��x_NU�aY�����{��8ܴv�)3�o�wZڂ�Ū�:?��ޓ_A��$u��� A�$f�d�!�^q���3���6�J���؇��Qj��!�C�-_�Z.�)�+�s����a@n�s����ۙU�OP9e���a��1z�q�^�6ҨAr���F�`�x����q���h��I>{\b�3K�{�֡�e�'�T��hVf��N��?��㹖�1�Dͳ��@8i��z
����G_��q,�����#��vᛞ��w'���L[���`���!��7V��ɕY�J��4���W-�/�1{26���e[�`Y���+јᛠ�DԳ�*v����f�,K��������� F�6'�4����;���,"�
�_��(p��J����{r���Gf�����M���b �
'�V-t��(���佷�r�|Ƚ6�f{ֲŉa��Lfyϴ��u��P��Hd<��1��Y\0$BdK��)#��x{`�6i� ֖o��G����H�M��&�r�j��Be=����!���/�	aw�q4��n��%eP�G���N+�j�vy���>v�þ;'B��=��ɴO�ha7/�n��W��lU�y�IOc���{X�9���W�.;ջ5�^J�"r��f�?��9���T�C�)EO�W�,����I%آJp/���Z�Z��}�Q���W�@!�����Ӝ���Xc}���'GR3�)IÜ�s����1q�0V�����|Ɣ�C0�-�͹c�ě�e�GM����%�4+�Pb:�UA.z������$�E��Wb,�a*�e��ѩ��b�P[x�:�2��4�c8��X`�ZDD�u��6���av�=w���D"Z���c�Hs0��]C�5�IS��*�,�9�D?y�/����6�&O���$-�3�Ι��\c�����D��w/��Ƈ��m����������&h܍C��e�C.?�v��4�@+�@�JEh�m��1YM����x���٫�דz1� g�w��f��e����� ��#�JVl
Ua��>�f@�qޗ����1�ݑ�9k4���M,=�v���w�D𗳰�c麶PF2�v�e��R���������Vp	��P\Q�F�͆�@x���)����)¤fı*�*�n��v^3��87���9.@3	G�H����u�����b��< �>�&��Q����UKR��W����x�x��$ɏ�uo,%T�ؗ��^�N��x���r��o���'<�XH���2�k��\M�s
ح�^�җ��I�XH��������sTh�Q �&O��ي1,y�ee��M�b������\�9>�t��;�;�Hk��ir�4��v�U?���6ĳ]�ӛ�?��6B��*���(J����==�ie�9��$y���k���HH=A��)/�q�=�k�5�Ʉ)e�Y������P�,8�����D�e- ��U7d>'m�,~��as����X��$�-�t�c3%�k�r��~�"���Q���P�OY.��|ծ�>o��[DH/�r��| �y˓h[�?3�-�i�in3y��Y[���wnR֑��4�u/qo�/&���7��:�<zQ���eAE�W������CA�r�ͣ���s�KI����9EUup҂͡s��J�wY�w�Z�J��:�'C���ۆ�x}��Qܖy0�Jp�� \KC��_��3|(��ggQ�N�noʧ.����Z���m{�(.��;�{�#���ZG�z\j����P�y�1�ӥ�����x-$���5��(-�����{�ć�J_#�L���S�!�D>��� �taR�M��]�G�S��b��T����̍�y���|�r�㫲��E� �,�+�.�+OW����A��Ƀ��p��ܐ8Lmg0xh}�l$�	���<Ha;;͏���s�0a����V�� ��۷��Bx�]�3�=���c���f�%9g��Z�X܏�r>�B(��~ 9��Nrw�	
�Ev/�;`$�.�8��g*�d�/�C��WN�K{c��<�Ƣ���O�I�6~� ��0&l1:�nWR���tt�&S���6i�iV,3@m�'j_�N�c���[8��_"������Ą��u���f$����%�o>e�W8g?N�d���̎jW�8��Gr6:p��[i�	�c���S����H��S��{�׵����4��A(�[��$Vخ��m���$>��M�����3ά�"u�������*<N$W�r֫��P?Z+1����vl^7ȵ��2J�6?�ku�3@����RR�:��^`��+g�!齙$�B�ד֨����(�k����ݖ��H	k� ����ߺ�i���Rݸ�5A��l�iX�����ܟ���rv�a�mJ������#%�#F}Rl�8 
$X���b�=�1�=s�W��v@��<~�e�D���6�N��u���4��C x}L������đGZ�o�/�`�g�D�*�}��Fr� �7#�b��d��)<���.�DJ>IC!q�?Vd�Ԭ�"��m5��9�E�S�+ #�J_5rfr�ɀ�c�䶩�}�R�<j��|�1��#�.�����7;A�\�׋����-Z޽ �$F�g��u��ie/����H�T��X�zdu<�o������p��I���X>_[*��"=�!�Q搆f�Yv{߫Ӫ�B(���sǓ�A��J����#2Db��vtW����x$�go�iÃ�l����R~+�N�_��F��*�.5>�=��Ȅ�f�����P@ǲ����'��䟁p�2������k!��^Ȼr1�K҃M��
�P��Ó����Hg,x���|~ 
3��B��]��}�LcnD�I "���/t�7�&�׭�-f.� qL�ͣ���=)�&7����Ŵ�@v}�6����p�^�Ls�B�����i�zֹJ%��� �qr�ޗk$o97��%GΪ
.� �ގ���]J�>��by������@㦹���U��j?{�8��eds���$���6�ĂQ;��g�2�:u<��A��;����B6#���$������놠�+!*��z?���h�#$�*�^hS�u�[�]�Y�4�x�92���Uy�}b|O^~�������t��KY��OƛJ@�'���T=�\Ϣ��!�5tQ�Hd���,�ѿ7Rӌ�nH��Q"��`
��sN3l�Iz��4���_S�(�.���P�LlI|��'��Xh��E��zG��O�J�~��i�5W���F�Zj�5�ؖ7��&g�b =�~M_�vxIPxĚĩ�/�I�F�������+���[�k���}ӂ��j9VԂ?�7�]�
Rl�����3�t�-��d�3X`~$U28-;�!=�xNn�)�5��0�#��l�<Bd�>�����BuꫝNI��������E�W�v-�%c�<e ���`�[l/�Um2�Rr����+�e��"�7���_���F�EPK���*��	� ��ʤ�hr;	�����#�3����b^0a�v�����H1��wm�>+�P�(M�(y�L����TƁ��Μ�ΒNU��C����Mo���@��-8�IJ�\�h����5��*Н�/,�����k�WkQA��9�7��;y(�E�vED���۱@K���߈`�F ��v�?�� ��B\��ug-�7��F��S��K'��c0��<`�j"��B]2mgw��B��"���ڏ¯C�}�s��u���[���L��M��Y��'�;E�Qg��9��G�+�lP���t��΢ᑫ���h��i��퐜��F�:��f?5|�Ë�
�|����@6/��3���i�8e�z3�T��~!�"2(֓�7�������nu��X]u��/R��h�8#�U�ڠW��#u��=��L0C������0�����y����d�m��yS��C}s��cG0 �1���A+�"�	\���w{!wF��5Û�;���njB�q���N?�?d��V�
���
���tÒ1�~X2�&���q8�,Xz���s���{��J�I��Q����0�^)��4���+�XMo�ƀ�8Lj��IB]T>����;�~H���!�;Jd�$M~F����;K���M}
|m�_�A�B�pR�T���v�K���(�N:���o" �<U;��86��|�,[c���r��*M�Ьp�sŀ�4s�H���R�Z��7�su��]�$=\��e\Q��\��v�B��|�Y��Aћ�r��Ia�H�T<�=v��ې��՗�7nA�?���:B����5���n��>Ny�a��i�L�Y,W�y����X�K�|��������c�;��<(�
�p�~��"Y��T�g��"���֨R�n�P�M��̹6
��.J%���,�ο���wC;g��"��s�c571'[�4��"��_UE���j����F�B��9uT�$T*�5E�1���� ���e\�<&N����rl��xa[p��_�L����M��n�5��<�=��y�"� 쾸9�oU��*�{%� r�B��t�GM�$�KX����4�:��s��2�R��a����$��j�̊DVdb+�U�)�<��˞��8P�^�~����W��dǖ��]�L�%�ޟ��ªz���Ln���89;���B��_���洯x�:{�s�0]j��'���{���&쵣�7?@�g'5��6��7�PW��h�~JU�����u��IjP�#��V=`n����Q��4���}Xn���c"@�7��2���	翏�G�w�\8�� >��`�T��W���&����tۜ�1�cj�1���/�W'ȄI;������I�~ X`�����}	�E��ӊ�z���sL���rs��\K����>|X3��ypT�Q]h��b0�E�x���vc�������H��@�l�A-:_����c��) ��#k,#��+�,��\���9����KO8z��.1�s�LF��c?;d�@S�͙2����/���!�o՞?߼�3��\QI�v
�^*)�^ւݯ#�)�I���e��6B�kVo2àlooLi�罻�I+0PTվ�_�i0�8Yzj �!��U�X�_��'�U��[�nW����.���K��Fd�����P���ÎbOe��$�JiB?g�|%��ǻ�#8度����RS���N�<�W��(Oq����ڀ�&?`��EFj�}��|�8� !��<���.N��0I�a��B3�!GC��V�r`NT�'�)`����15��,��5�%��i������:���n�LBp��N��Ycv�okuB����u&�ܬ��,��\u?*��?O!���îѤ^MY
��i66kb]U>k�A�p����m�K�(zG$�9�s��E�)����:2�m��JR��2�ph�!h�n�r�l��n�:�t��鰺�<���㗖���Qq'�Ϻ�{�`�//��9�;�k���[�MU��p0�N����M�y���0��z] #����;���rk�4x������x��4	/�GKSVP)�	�S\_�`��VV����_�4]K���=�T�a[�KO!��J� �q���Y b}�� pEN�v����L�\T�U��N���.\�s�tg7�~aF 20)��7��ǌ��չ��>����e���*��KՔ���=l%��3B�:ꏄ��,]������$x�'"��q�Z��UD��	�w����hSL��f�U-=�\���e�L|\�㡠�����8J�U.��|�5�d�~*$��{p���L�I /Z�"�>��k����JB���8�x6��'�<�z�6z�	�Vsa��B��}����&���@�}n-�,��ǩ���q"T8^�J;2p`��8]��c,�Q�g>�G����z�����9<{W�c���PN��b��uV?���'�ez����2�W��;�2X�T��˖=�������NQ?
�m����èC���"�lZ1=x����3��8Y�>a�C �V:����]�_����&�0�HĶ��J���������O��K�`O�.D�A�#������z����6�2�7�����X�zӴÄ!���c�b����ɍx�|r�X\{����!(�#0��s ��'F��?����⡔&��i����O{��)��.�a��˪�G��8yQ T(
���LEP�Puø�������Q��%� �{c�����X�o/���$>�ri
�ۙ]
���5y�{iiЏ0�z�V���3�g�e\��`�n3��qӈ_�>�5��3�~�S���|���P�Un�=V,��x��V�;H��0�2:��9Ph���o䳯 ����G��ʹj�\őTg��-P�ZL���oОp�j_V�VӷyQ�[����������(��"[������d]��&��U`L�`8	;d��D�E�r���j}_��	���ZD8Dyx�xύ�On�=����=.��u���̙�0@w,��גƹ�[w;/�� a>B&a��$������M��F�>4�o���l�e��}[0�������P<j��ͪ~�f	�m��+�g�3t�۵�jb���5A�d�:h���z����F�����e��6��p������Z�H������.KDt��b0.��4�/���Z����g[&|�|�ɳ �Q���9j�!�	`�˹�g�D.<ըF/�n�.��y��Cޘ4��]�܏�������~������뉱����=��;M�����]�3U5�%By��|�5y������UK��œ$a�-����*�&;V1�Ȟ�q�(��8��ŧ��!?p�ع,�q֍��M�`�x/Ӗ�2;�{���f���E!���ȳ�p��YP�4e��uO�jy�v�f�$Vp��-E�ڞ�fa~i���~u��p_�夲�g撝�,c�2'��Q,)*ݔ�_�FɟW��M���74���1-��q`�:B��T}��L6M�<4yǰ���8z��T|l'���D��G�F|Ds&��2�Gۨ�� "h\� $n	����4"ml��F�ّ|����"_ヲ��<��$g�(D\�"��\Ӟ��I�?0����r�f
X�i\&��O�����|�*�'Kz�G`<��\S)��{|����n\
�$	�Uېop���S
.(ȁ(e�~��۠A��o�VŁ`7K���n�·�5>�_���=���QRe�A|]ςi4*���� ��"�62�ژ���['ʻP�Y�Ǥ�ۡhO�r�����lX��*I�4�� ʨwN�΂4ٓ@��3ElͳI�=M���^Qעqj�;b���4���b� �z/ ]r�oDId�1����Q���gl!��'ƽׂ7������V�Ő�� Z�Z0��ն�ʧ�y�`9J�Ԁ��S����4jvy�Uͥ	16T)G0�ѣ
��3! c+Y�z����1�oZ�qF��Z����Ren�j�*��ؕ*��a�`���#k��]�kb���d�Zo�h`�Ϸ����eh�;G�`HQ�X��2��UU���'H)���.�� '�y�h^	4�҇?� ǭ�}�Z�� ��8�L�rL~�#0�JK�8���G�`S��Za�`���О�x�]{�V��)>q֐����v�T��9H�x�s$&�	����pb�:����v��j�s����L��������`7Y�"w��8�ؐ��U�˂�.��kW�q5�����e�QkM��P[v[,���Z��Li�Y`��cO�eW_���d�*��众�}!�1���5+g��(����)��^�P5v���c��D��;ke.�7��fi�\�xrY����Yr�{� b�E�(#=	B�<F�P>%b+ F�}M�-#ő��ӏ�[�]I����e2�O�J�w���F=��'R����͟��
e~4�M��I>/�0]�T��"(�rV�0��\(w�B(�͢��%�6#w�!�z��:�,��1U�;r�N�cyɏ*c��Y��O�����u<���n�>�f,pi�7)�!�Or6\�I�!��H6�lv�m�H���Ю��C�@�ͣP�������m�h��X������= q>�0O�g2H�Ϙ�F\��뷽��E��l���s�j�f6ropU%wF-j*!�f�6���ڱ:G
�A������AY��ù��l�9l�Ԅs�L%��y���^q�g �.���8Mo
��Lѣ�J^��s��۹\uE��w"J`�i�J)[-OB�M�n#݈�d�Q��6����Q��`�l�>�g���;b��!���s���{GV����[:'�@=8�C&���7�_�[����p���uFNng�� {���~�@DX;$?j?�N��K��W��D>C!ȃ������/Eܯ2Z��L�~w���	FL_-�#e�
��dP�Ж(k�`�\�e�?+o���*�f!UzhEOy[�9�xѵ��9����.S���ِ�`W<��qqE"r��� ����٨�9:1<�.��D�C��j�<o
9qTK�` ��*�{E� ���>��D�NX��Y�����_ �lww���p��¯m�A7���y�o4d��9:t��5&D��҉��qR<���XoOLZ6RDX^l��gg��k��H��y���+�HIcUo��D�j�/�IF3�Z�A��+�����y@No�0?G	�\ٽ�gb.����i�$��.�������yⲟ}���.U��^]�@��=_E��CV� �T���5�>_v�@��Y��z@b��uO�Ff�%���~�"fs�a�$�rҐq��"�� �e�D���m*{�pl)��v�m1!(D�?�'�ҷ+�)3��)�B��@��q��+��B�w���2Um7��H�Z��7���1�O����m-����1�e��"i����s9j��0����(JQ�}T���"M�L�Q�騽��n��%f�!"V�b�V/���"��Ylώ��I����|5jR:�[/��fcs�!�l=��vH�Iψ\�}OjEX�^�(:���+�$�֤�>��v��gn>o�͗7�kN�4�h����Q�D 5K�o��tT��z޻w��Z����7�Ը�H�C>�w�g��5���.�̭i��6�� ��|�z�i>�$Jw�����@8�drAc���#���� .+�8T�I`73����}��泲T$�����=�QS�>cǼ
�Y����n�?��F ~j_��.�q�Ki�M��a�Z6H��1��L�ܱ�oys��=|��a�-�^-�:��?'�Z� ��� �J�<Q҅�;�+����N��g,཰�ZNV��}932y�0Tͦ�l��_R�\툈�>��F8ŒK>��w*k��Ew��XZ��ͽ��w�I3׎���F^��M�τ��X߰����|�z确�
X!�G�/l�J�M��2��n�S�����.�ί["����C\a�#3��b%�\��I˘�ߦ:e��-~�9��vo���Jo�3��<D��渊�'����5߼�s[�`���v��_c������R6N������p�&(��S��(K�1��=
F)���`Ա���G����>��c8&�xԸ���[����v#�����a�0/�P��G.�"��2-|��k���^sl�X�9�C[�4�eM�a�-!�����Z�&�bƩ��P�fп'_��M*�~/�r$/ ���6t����^�	u��U�S��!�~�#,h��]�k^���ƞ"σ��aD�$ҍ,���!wh�0o�ld��T���E�em`�6�Ir�ӑPă$o����}�?F	�����7�+�����ܓp�z���y�8^c�䥰�Mq�Z��[ݗ%������)�ij�ij]3i��U5�1�,e�u�,1��s$v����n�7��֒���j/u�mƌ�<^H�ɲ'OLTZ��l����W\��/ָu�[-�+�.x���>t��W ���1�"���J�J��sZ�G%�I����"��ҫ9p��"� "����{d s��=�I	�p��"� 抅Eo�ֻ�gC�<��=u��	�;'�N8hǬ�T�w��6���2̦~�[�,���ɊC�.Y�PF� LNO	��2������z9�%\8�ţ^r!��k:�i�I!ˉQ�:�j߫~�ꀈr�5`u�Hh�p��͘�{�n�u��ksO�c�Ϳ�P:(��]�rw��'1SǐԨ����,TԔ�����}�}����>�&�ɷ3xb�\j�."�J�ӰL�*��Ac��l�t�1�j��3�NP��0���S#�l}`��Y���,��p$�L>��ޗ[�U����cI��{����6�$��
Z��N:�th=d"��Gȇź*��u�t�4�G��_o�~�`���'�0�0|��ʁjx�4���o6R�A]߮fǖ��>��K^��goYDD�ٻ侸g�F�-�p�$E|�	�)Y@;Կ�8�������~�A H��l�w��d(c�Y�3�vH�|	<� ����{G�/�|(J�fOú�]h��]G�	��ѿ�8�����ţ�@�jy❘[�	�C�<l�4�/�]B��:%��I}�16-LU�� �oo�l������������Y�}�k�P�^�����M�=u�<%=D!����d<)�M��)ء�du��K��?N��T��*é�V?K�}c���	�5B���[�k4�����>M�151����0m���c�A/�-s8K0�	F���j�>���X�-ɠ���
�2֬-�u���?�*�?�
N�Ɖ���^��u(	�~{���`�t�ʈZ9PRۜ��L2�Ki�SN<(����[���o�¹��c��̃�zZ)���ص;�����O� G/ix�B�PFe��?��
[�rs4���fgJrhOWw-��3j�\y��H�D4�@/޳9�pJ�֭�O�dQK�ez8\<�V���#^mΏ4$��5j�׿�MBN7�.�6_-��Tn��A���!�9
N���ؖ����"Z]#��e���Zdy�K��`��GC����: V��1�˿�^�+����q�����V"���3���ߦ��$���^�:��ekS����)�ٿ��<~)�mPM�G��G��(Y�.�V&�Ԁ��T#Pz��O����D\⨀���R������hW��ܘH�,����Yp0M1���'�����u<��pA�E/Q�F��� x��=�� �jzKF窴��J!ʎ�S��-�Ap���2�ɑ	�������b|�}�<�;�.�ކ���(��=T��Ev�7U�8<<��BڽP��r�1�8υڗ4������eAŝh�G���k�,�~�+�9���4�	p�sJ&/�����~I
�gLF���#���\�wG\{G&hʫ��x�wBEQ!p�:�Q�
H����;��2t^��'ӫ:�s���P����*�M�}�Ȏ��§^��2�}Cx,���hE�䣆�]�rE5;~mv�#����3���n	�)�����|�{� �J���G����RuBp�x���(��4�z=�O����*D�+�ѭ+j,&Ў	�+���Mt�q�I3� ���\��е�9�گ+zf�Y��F�$�i��`��������f�E+���en_�W��_�F�3�	�$����6k>a�X����	�W�l�����#�� M���*�ٔ�d�1cO���A�b���`�\�hz��9~�����.!0����(��-�ҕ���ߦ�@�-���H��T�,�{�r�����=�2V	?������n���m0��m��������t*�;�۩vz��S�&f�^�v��,)����&�k愈°�	T�i��M��Ӆ��cA�(ʇg��[����V��z)W�PU��\�o�
���0f�S;{��1ˀb&&���UoQ%�q�'�T�g=7��a!仜�� +9�����=R�6L�ɵpG���K��߯�H:?:o�N�d�
}�K���3�Z��8�u=p-�s�2mq@��wW�n���5^�ۧH�������!IП����ҖT�p3~ۖ΅�����\bBE-�8�t�ѕ�b�Au��-ĳ����@��:@�}�x�'݆V[�����Q�v �M�Hr\�ІgE�
u}�K�@���|��%s��ٹ�t��JoQ,�9�0�+�F�R����"}�Om�ۗ����.��'�pګ���z�MT��RY��Bl�S`����ߕ�1�D�ɉ��c'�=qG^ggm	-E:��������8`t�iUH�F��~,�Ob��96�;�17eZ���8��d�߭���!���ɖ&�l����U��x<9�G9�<,�Yc�fY�K�sZӊ��/,�ص�����_�B�>��(6(��8,8�y��U��f׸��u^���u� ��b9�%x	�|�$��F�Mb9_��ڻ��C,W�P�.$\��Ŭ�)x���R�"r��ۍt�L�5s�&Y�X�x��:���R�N��A&������ �+��dg�4�B��@�[��Q�#�XڃZh}��/�z�?ыa�����5�/�O���]��>ڴ1֖4��n5;W����(ē:@)%T�z�V��D�;Ԉ�3P��3ƔQ�j� /R��~t�Wc_Ƹ,R�V��(�	WM�m�W�MP|3�i��\R��N��~��;q�p
c`�����H��|;vꤔ�R��엸��UM�\d�ʭ����ͽ�<���hu���񏤳[xIjw�_,恹l����B�8͡���֣�B=Un���뭔)�Tؤ*·z5r; }�q��>���D�B�q$;,�%�����# ��,�ںu�v��%Yz+V@�64���z�{\/f�?	�l���5q*�E,Xe��F�1�{9E��f�{���1]Y}��ҧ<Fl왅�V��x������ɼ�k�Z6��p�5�w�k���(�@�Q8����\cI'S�V����lz�>le� ���(�W�� <��<$W����7/�l�s�P4[��!̓E>=���H��ȥ����������1M֚@n�2@���o���U�F�c00��<��Ot�{�ް[�k䙀������v��U�L�o}E�L�J�i��h�^��N��}�_����ܣȚ,�WF<�?M�	����l���c|�E��[��������-����vb��颡�ρ��5��L/�{��?F��̾^�\8R��	r��X�����ބ��}��r�HWQ�DO�����"��U_��w_����*�7�f�^����Y](3�����" Z�����S���:N������G����g����(�D9a�o��͎ݽ�� Qɓd*�h��09�*e�?2��IC�Z�׋8��Jk��ŀ�/,^LOÉ�v����y���k���S��px�����j	$C��� ؎���ؙ��i�3��]&r��t~	��r5���}<u#��A�Jڎ�7���q�Q.��N{�;uW�1-�B_&�W�$�1j��8W{!��k����#IE�suW����h;�H����	�<�����"9��EAv��?�%P!yҥÔ%i
:4��xk�2QY��$��:ݑ��n�1p��A�̔$�������,t7�r�Ru�m������9ˑ��	��
CT�`p8�nD���[�7w��R\��qQ]���>��hƁ�������f!�����ϊHI�x�)ci�s@�J3��ʒ�2�v�@c��u���_ ʨy��"HI���|@���$��b�|V8�����
��c!.׹�ej�Ѷg�9=9�%�j��,��cx�d^�o]3�X��)�`������(/�=�5�� S��)j��F6��A3���9�E=��}��L���YP��.)��s�[��Jķ1!	jM�=jzQl/�r�RCjX]�8��/�ξz��㓬��j�RA��2/J㢦R(����0�l����a�<��Q����m��>�%tB�^~M�cJ��0uG7�AG:\�����#ndv��F��ӏ�e�ې���&��٦U����diD���R�Xw]�M��A���[� ��*�}����:�rp^wfl7)��(zT��j:�����ji?rQ���^�րCۏѱ�%s�z�zz��M�ۀ$KX�9=_U���1qg\"��h]���'bf~�4n�H9C��?����f|X;�"�zA�ʖk~j�ו#���O9���==}q����7��s'����I��wA�ľ{���PW�����w<�X�G4�Ԋ[j�F=*���]%륓�==}|�G�(z@-I0��}(��K��ZS�7��PNJS��F�fv�1�π��)���+��{� �x{H��2��%
侠����>:*�S���"y����l��W	E�1~���y縐8���o~p1(o��`�w_����L���h�"��߿������_�� "��͞��s�g�����@8�#�>��
�����R�>o�)�<{�?C�jMqme0|�ʨ1@��(@��30��\nvn�
��ˁ��,�&�g����RCS��;��\�s"�[_{�`X�?a��:�!�{��*����N��� �3A��,�Z4�5nh"HS)�v�=Y��9#.5ܻ��v~�bh��V���\��A�|��
���V8%��N�`46�X�E��|�z�K2�6q�B<�|�i��.�P���j�k�]�T3ť"Ȧ��D�~r[bߤ���#X�R޺}���V/9(.�;T��n���Īw�x�6�ҧ�C���Y��Y@�~DVފI�~�_�c��'��Fk��}��9�T��|���~E�[�-y	1���.�BCǒ-���Áp���F������Ġ"��8���h�e��C�;H�@�5O����]��hU����3?n�Ih�]�X���sOf�85��W�q��� �ʭ*���ͷ�����ޘVt�T/��H|X[��\�f�lN�I��<�ITO���7%*��%���S��c�?���'ur��k��׎4�n-�8�;�'�[�!�����ـDRO�R� �dx\��C�������j�u�Oflv9}"�h��d�����"���6.�tj�##޿\wH��#�tH���Z������.a�W֮�5B�r�|�B+��C��"�ӱ���ò������X���x(2u�;���x�}���M��O� �sĹY���D�宯�yT���l�F��%�?��:�+�Yy݅�AZ[�0�;��q�Hz�#�Fh5��ʣS�Ibb����=�����	ވW�0'�Bٕ$'&(`n�Q�wc
kWJ}3Α��������GF��8,�i:���	u)�9h�V�����C�>%w�U�n��l�vcȣ�H���.},pN]e�BCc]]�-��[���Y�����g���4�%�){�/��cI�w�[��=3����m�c���7�HPVt��bJ���C'��6�#�x���܋	����H��Ιo�BR3���� ������i�m)^4 N�g<аS�}uӜ�g�{e��m�
ǭZF��@Bz�E�cQ2���: bi�H��s�A�ۧE�,6��-o���W16�#{�>#�z�q���$*7(@�pΜ��ì}�J����Y�]��_�p���U�̨у��2l�����F��WKs�A�%���ff���廯�+Tݽ��E �x_TcZ�w��)����uߞ7�r�$772U
�N�fi���ٺ`�!����e��������8�aU�B7�mc��l������4L���/?{�A.���� ��
�� ��9�ْ)f��QA��0ƾrw��݄��3�����<:TiȂ�0 �����ÔK�;��}��ɟ���\|!�:�N�����')W�zT� 9�A�U��P��u�=�K0؏l�):BW��W�|����dog}Pl�����bN��Ow����9�l���,.�%�)��ڥ��NX����֑/�Oֻ�K��niΩ�	x~[Ene��x���Y�좹������PO ��YӰ��By-��Z��6)r��]EYo^�G������[���&ћ��{K�SK�s�����v�3��S	��8	��s7���n�wF_c�	3]����Lp�o\�g����8�ޢ�W�h܅�=3�`>OHƅ���6�~� �t8��%M�h�"���Ѣq�k��\��:<z�^�3��}�K;�Mc�ԁ̰�O��Yx�<Р��P&Ԡ��U#[�V�$�Y˄V�'�6wbj��F�e#���z"�9��o4B'��H!�����[ǯ��5�����ogװ75���QĒJ0W �ͣ������˻^p*��6���2�̗��ۨ]�H���j�>ݼ�B�H�~w[��o���Q�y"FuN$Wa}�hD:��jx�ȰD��6�R�fyY4wP�o[Ǡl�L�zP2���~e��g��y�'#����Y��\E%�ʨ��f���,̯�Q��끤ֺ�*��(z�9f��2@㠳O�拠��~�e��&�+S�"*���x��iG�FN�\�{/�3�|������H�2��Y܀���is�I�Iޙ�P�&��'��^�)=�''�|�]"���S���"�g��B2i�`;5�8��l,��:Y������ pͼ�%�{ %IB%N��e	�#QZ[���m�P�x*��M�P,�J����K����1����ŏd~����m-��W���	@*�G	h��L�`� Ɨ���'@�����C��c�=�Q�hn��l���ri�@��N�C���B_������O��d�'o�n��7_t�q�d���h&}]:�t5��-�%v�{X�xDv��p�l%/��"v�Jہ��\������eD��s�z����Z������ ���T�n��k�^o��/ �g�O�?+����0���D���+=Ǩ������dƖt�Ѹ/���<��\z�?�#ښC%jM�o�_���pz s��&_?u���&jr�-�b���R鴟bix,w)'��U�����O��gu 8�K��ʿɩXAK���KR��@As���C�+������<`�䂉�ulw�>��y h��p�>ڇh�
��<������a1k�.�l�Y3�G�xG��|dl
3�A�A�ջ�J��}?9B�&�y�:&/)?��較n[(����s����(c����s}�t�p@��d����	����E��L\NX~1@�����yvx�6G��:D�"��{��Q %�,"@��1����9v}���~`�~ RhQiz?}��r��%+�]�� �X��s���Sja�˵UO�$��r����5O�m<ϊ���
)B"M�ZU5��X���IYR��9��y�;*��zJԦ�u��s������0Z��`��~�g�uV����yj�e�h�7�E�e�)J��-N��Y�`��#	��_e���ū���pZ�pZ�K��6	$�{��kw�v�)�~t�OWD�	�5jq3�!H�y����D���Z��̤݊��H.��	�&[+ggL�|�/L�|�`c��I�J]^��xF���l���.u�ٜ� Ԭs��2�SZs�xƒ`B\�4��0<ru�l9���
Z�=RG�f��uGW%�k`x�E�.�J��u:(�g���`���$Y��i����8ȖU��wu����X�4��ɀ�W7I_»[`���s`g7����N4�?O�S/��M""�9���'Fܵ�uR�9�v���]����W-�YJ/x-_y�����b_~;F�Y�{<�̬���P;�
s|�%�&�{�Oh��s0>Z�6�Xx���N(��H�|'ڔvpG���0C����2�=D���]����Ř���,E62@���^�� �0[]r����A\�S��`[u)�rW�85���6��԰�"<cd�G%�ƨt���a\��n���E\u�;�2[g��Խ/w\����`P��f,Չ>4��^�ل��A2�@�M.�V+r�=���eGr�b��ڭsL>�HR�H��[ě�#4��#�ݩŅ~�Ǚ�}B��� ŴjKZ�<�|K�rz��#�������i;�|��cO�>ؙ� �.� ���c{�04~��B>f�l���r� BD[�!�d�?���@�/b	1̠քO��l��rN�t��>�qo|��`i]g�2+ۯxH��cu=	`�-������A��¾��[��V[�8�����Xx�q����Y�}nDo�C.�z��
�!�릁2I�x�)�&����{�+��`5�<a(��n�m���|����7�&�y��<��/���v�T�k=��<di���e���$	��У죜8s��A*��gUSA�/||��ui]�3�IF@6�h�q��[�G�.k��}�Jǟx�4���ua�XI���#0�s��^���{��f��k�D�������U?��5���4�g���c����[��h�	I�څHG��J���ȚBɥ~Kk�}.���D-6����>�p���m�N�z�	P�I�m�7_�[=C�D���k�C�e ��<�7埫�4� vW�8,Jȶ��vr�b���_W3�n�0x�n���9_�uK&��W�r𸐥�43�b�ռM���l(0G+aHs��|���ދ:�7$<z�-d����g�m�-&���C�^�i�z�Q��������������K���e�|��4l3��&҂��}4;�Pf0*[���4�Jˣ\B�N2��h��vR�-M��Խ����y�\�t۠���X C�{��c=�۵c.?P@�eF۝���g"�nV2�]����k�b�c�W��?C�����'lOhSQ��i�s#5�p������\��L2��ylz��5x:��R�$���/��]�N��-a�kΐ��iBP���r�5dkKv�$�#��=Kr�T�fE��9E�%r��O@�B�~�K�In�@#��|����l�'<.t���30␩�3���3�Ϗ���'C���s�|*4=���:K���BM���ߺ��/yNY�D�i���@M�@|M�`?-�
$�Y�c,w[�H�_�t�%&����%oC��+�\M��	��Qo��}Ҁ��S���ߓ$l����`��z�3�ߝ�;�1�d�l���2�@"���$��ߺb�I��i�D�*PɠPa|��v/���~g�t o�o:(�s8�tάk���N�T��sЀ�� f�$H�A��*��h$LLe��ᦗ?�&��S��cS�{�'�)�ī�M�P�nf�L�;�~����-���_�ԇ�60�GI~���À3!���Y��ѐ�6��������w�2.}����7�DSpCu.i�������_�e-����!XήX*:�(���۴Y�:�p���?F��E��;2�R��=Ev�[��-�s3�1z/u�v;��=�������B�3�,<�̵Wn綡���p/��N8B�C����r�t���ʏ��[��K��e8��v'7��e�� �G�wE�l��Z��Wz�'�w��V����� �Ri�����*�dC��,�oJs���t��~��	W˂�<��B�%����Iu~��n:Мh���É�	?������B�8�>/j����S�'d��(D������_t��vf�G�t��m.}�:����zau��Ԭ���������p���ɇ'��go� �����yukwn���L�cr�/��65~����'�w������6��.�J�]n=w
?t����7EA�⟖z����
T�����(Gx�l�U�����+Tu�]���TH���木+'�����w��Tad�:�y:$w: o`
�Ա��|Ho�{���C�P���B��P��N�kX�da��,̶_����@�9^�¢_G֯H�Al�����Ɵ��Zc�pB:J�����2�+C
᨞s����7��?�Q4�J�6q,W_��j�\)��*�����T�[F��[4rx5��U�cvR5�r��f���%L�['�y��k#��"��=QR;�;.���v-�� )�m���`�L�-Mn�,i��>VJ)��_�,�,��܉���/E�����-���9�_�圗T�6VTf*V���,��3З�(5�P;��Z����!^�}�6nK6��l�\Ys&<��/�č@oh�
{��.p�gIQ}��yV�Kg��$x�sD� 7�����Ś���'`#s�c#hx!E��n���v������i��d��+۶w).��l�V��}�h P�<����V#ɯ�Vl%-�<	���M��2�3��'�)��3����b!�s*��U# ��T���A�y�DѼP��!�P��QR��Mo�z��k���<ռGg��Ӂ���a�F��e� �XG`��F�
��j�C���*ۂd))|ZfK䧜^�^�߼���HJ ǵ�>��~��.��Z�F�h�>FY��v#�x�py�m!�>�Hc��K��d�d[�r܍{�������ޢ;�׃̵1�d���,|<�Ri{�}���-]^�����Բ4:����P�Bm����P��n��nA�8Ϫ����4��R�F.�ҍ�K��{�Ira�3�9��TM=�`"9�V���I�{e؉��τϿ��v��D�YC&�S���l����ߕ����{��Ki�6��k���n����a��=}�O�_�|e�>��'�I�e!1*�d0������k�6�XmuJԕ��X '�=@uC
�(<X�a���&e���_���O��C�����l�5�C\37�Sr�/%@~�	෢���%$�ȶLC�9��0�����sI�ץX1�"�H3���%�a�>o�c�lni�=�Δ��(Rn+c����/t�7�]U��N��d�j�b��_<����s������`��8'|�x!�H�K~��&S8�;b��%��BA.ls�NV�x�}0���v��v���q^R�5ŕ��P�MK-f�j4��s�J?�Q�!zH��9��t��d�M�'>p��x����S�:4g]q���h�b=��w��4�xP�\Kjڽ�V�s,ط��-�\cJ-@"�j�z� N��������
$&��Q>��"�@�FUy<v�pcT��* @5?Ҩ��5����ƴ��#\��^�H�l�nP?y5;>#�w��V�i�X<D5��Q�>
��Ԡ���5�J��ʸd��������/� [ABp�~{�����&���u1f{
Po�LF��[�w����`�����x��v�i��t���+"�3�@�U����I�#ZTJ�ܓ���=J���YJa���c��8?�������t�P� +��p�V�Z��!���X|U �.&T	��O�^��	i6:��������;�0D^�mY߳��`J��w͕0���W�ɮ~t+6�@�`��>�:gqf��A�d�O4���.at_E�G�3܍�f�\�X]b�7r�������}P ��P��i7QB��MrQ���I��뇫�1�U���g��40��S�� Z\��=�����:��k���ǰn�Kk����`mߔ�Љ��.��rcC�w�lO���<��wj|��+r�⦱�`�}Kߤjr
�³ȉg"U�|������U�q�Y/��c����)P�͝cB_�<��IhѶ���|1ݛuw	����#N����h������*Ŗ�	N!�Σ��?��
1)N6��Eo�۱㏧�@���T���Tn�(m����������<j�'�*��O��khM��{�F'����҂�Ӧ��@�D��1	J
.Q�G��x�V�I{�7�O{rXN�Nc)��mϯ���S�DE�Á�[<�2UKq��@��G�G
!3�^��e_�{��@K���)i���54C�k��dq��P*����;�М�cd6���Tex���vo�8w�i@X���oQ�;���2�9�A��<�*��c���bxH�Gn�h�/#O�gG����P9�IWC��{��"��]޳�������I������}��������gZv�/�1Ʀ�x�ㇻ�����{~�yg�dԒ�cq�|�o�-gDC#pz ����L4� 1kzh�4�Gw<�C�6�s��:a\���-��5!|�:��Ơ��"dUnn�̩�=[�����p�J��S�;]QP�2R7lD�Wk5L}a&��eZ�f��ޚ�>�(Gk+r� q��ɉz����Z�
\�uu�W��4�)X�O��A��Vz����Q9������S<���7�}�?���fDP�p"����>�TS�N�s�8�H�d8�r� ���06�Y��������^"b�y�`dǁ�F:����2���x����I2��y�-��	Պs���tI{Cۙ:s�kV�a�T%9.{d����`EƸe���B��.b�i�h.,�9��\�%e�7\��t���L��~� |,�|lٚtQd�2+F�u]��v�0L�aV�&<)��|��� �� f����f�guw�h�ƿ�7_���$A�!=��J;�h�ROra�����s�U[V�^�z���
�V��όu��՛��ȅ�b��>S�g̳���î;2�}�"�����-�u��3�,����)��C�d���6��1>�P��^�.$1w�٨��u"��1�8w��e��#��Y'�&��e(�"KӚ�e���m�ۆ����ĊVv<f���C��y�Y9~���d'��IAupo�	O���eʆ�&��_L�g�뀬_I|��q��V�_/m�����l�jJ�����U�����28���_E���K!��ɶ64����A1�vNA�G�e�l��f�ήrbO���(�
}֏{�z��=��������<���
�7�beŏc�2<��Q��c{*N�J�@�1oÝ�wT]\�*����+9�&Y��a�׹ű؍.��P^�,Xt�Y��4(o�;z��8f�9 <���|�(!�e?�H�����H��_V�ƪ�X�m�>�ֹ� )l0v����t�;S�@6�:ތ�s�q��n������(���#��A�L��W�O�?#��K��}��Zя��׵��v�{�9M oV5v�X���{��*X�]`Kk��?����Ns�G!�:|��e��`�s���iaL�]Bn[k��l$l���ͤ^͎����啁��d�[��j�8�䳾m<�Xz���&n�mq�p(��n'��i�B��F6vyk��wJ��}�Ҽ�2я��u~��۬r���ڍKɂ�^^�#��9,�n7p `�K�j��/1p�`�G3��o�j��6�@OE�
�C�aa��r��������	ƴm���G/�g��}�`k��՝5�����{&�_:9��=m�%/q��/[Ӽ��;4[����n@�p�&H�kV���1�ϧZ��f�͙����ڨɘK ����E�4S�����)�Xm]�W͜��c�1K2Y��M6<6��(1Iv�ȝ�d�rf!��
>�,.���B�%�W� 3��yd%�.�r;�
K�?�(X�ǭ�Ym��v�� &��������E���� �n���
�G��ʲ�A_!�R�$�:n:AȢ�W�Hc�q�_�#��&����ډ�T�%�g�-�q?+-�R
�&�9�$X+<�o�V��eg
[4���|��FU�r&�����^T����������/�C�����zH{�����w!2�W��o�*�¨y���8�QҎzD�pAia����-��G��B�D��ª�I���K��[a�BI��}� y���R���H��8s�u)�ݷHDB>��;fh�-�i{����{��򜰌F����h7薒[� �8�8�W���I��k����2f�q='�G���p����q��BӋ�� |C��0��F��:TR#},��0�8ܲ��cMؑ��5L�����l/�~J���arI������РɈW|og8a'��Js�!�*"|�
�勸�x��\9��qU�G�&���j珞\Lq��j��8����=���u�z4_�%e?}ڒ��T?��)���
C�hB�/�]Ϳ��R�7G�vn-,���� �,Lw�F�7}a�>tkd���ڂ�m��LU�0�;Ay�ͱ�?�K!R�æSƠ�f�S�*�3:���$땤�\��<yFডA�1����"��*S_E-�H�l�mtp�uOv*rȮ3���ȴ�LL'��$�Sp��Ԫ\�,j"���o����?7ꑩh��6Re�ݤq(��+���śׅ�q*Y���b���?X�6�t��b�c����i&���"��O_)�>A_"<x�|
�Y7@��|L��린�y�غ��f���zň��N���yxs�Bˢj�ڹt/\�{�b�kd ��5���-�se�}a5BD�rn�0:zG�@	k/d�����[j�E�[+�e����:��R��8�{gv�� ��f`lq�����$�11�Kop	�C��ݛ�P*ū�Z;C�r	��<G��x�s�f��2��.�̜0�y�?����7k�p�Zh�.��^��R|��]`g̗ݑ�s�G!�G��v~�êTn��>��eT�O��ҝ���۬�(�x[	�'���,�`�CY�QƼ/��61�������-f��#M͙��XgRݚ��;�� E�h�8��N"h�	�$�$nC��An}@N�2�p;Cz�M^�-`H�pz)��+CW����It�TQ'���d]����'3=7��]�����.���йs�}�'؞{�[�<�F����u�q����x���@�)�̜�<f�zϋ�끭vi��N��˹,N|�f�%�R�v$�y�wT+�a�q1�D��^�Yi�]ỘNH�WB�ʾ9����i�7Oh0�5�}EJ?C�;ŏl�Z�)�}~^�n���5��hB��(��|��C��Q�o+���X*[���JR����)�	� ֭}I�H��ǰ<�7����_��Z�J�����K;�g{��Ȯ��	WB��wK����˭��/X�K(D����-}��C���zPI8p�H�0o.6s�s+m�a��xUbd�+�͸4�����ht`Fs�ZŲ� �?q�fO,Ϟ��M8Z�k�.A�^�?��- |�CR&�ۡ���s�aEnM�.@���'���j 	D9����ܠ�|�>$(�y{�W�:�D����m PFI�VD�҅j���_�J C�F�+�TKN�� �%r�T��y�[�;�*�&cq�_�'��՗7_�i��Cb� �9�"@� �p畢-�Ǥ��	�|��p��0ފ*����[�<�����0��ѽ�����e?����`T�dMỎ.T�����/
���,h���
���{D�:����ȻHH_��L��hc��}�8���E8(�GQo"1�b\���;j���OJ�i~T$(C=pc�����fc��d{9-�ͦJ�Į�=j��&���﵏
v�����*Ld�C63>y���/�l���D!��7�K���C� .W���J���Ϛ8p9��h$B���r�M��l�2�b��X����#�Ճɽ/�I�P���("��<錠�w��w�=Vpv�͍k�@�y�T�:��1/&�?��z���h}��~^���Dj�z�� ڌ��F��s~���OO��ϻ�\�QDi����� ����a}jm�n��]�z��"�%��w��c��v�!�M/�믮����{��y_���'��p_ّ�Eb�7�ٞN�`A��&x���*��4������8�6�uX�~��2��R����+Wk[Ax���A��A�sH����[k%�����?���<y�ţG��=ɗX�</�e����<��WN�j��(�M=����Q�9��gh�.�#���#��.w�C%�f��)� U��t+�=��CP4�&Y��1�w��Q;�
N}��'�ۛr�q�qTB8��A��Y��R�Y������NJ8
�:!�(PgㅉҴw�� i�&-��2�����L>)P��1'(�__��Q�����P��4}��a�������k�'�؇����˻T�X��:��z�yNg���]&8|�m�f\W���T�+�WQ�D�v�nT.�⠃��^W�y�7,���J���!�o���%úӬȐH�T��ܸ�{���g���OC?ɠ�wsݫ��R�ϪO�S/v���w���	.!������������r���	�F��Ͳ�:u-������[ڃ՟hE%b~=]i���6Gf9租y�(-LpG����"��
0���t�݅�%y�TW��k�nW�\0��NtM`S�Ǻ��r�m[���t"����0k��H�&*�z��r6��Q��;��g�B�F!e�<���_�ُ�6	����7mT� :8�&�n��NP��U�y[']&��a������r3���m�}&�߄�~�D�ó�],������hoC�7��ͮ��?j��c� &QI��	p����6h��ޗu���P��#� م�l�Ǿ}x�`,�W̡N5��#Dʱ���8Vɖ�6o2��G���z��.Z��4���n,��V��{O��?,���F<xo�k|S������ H��<|k�4���E�5qU��~�B�PȽ%I�	�w �8B31sfE#�C�\���?�wz����p�:�������I����`�B���F�s���d�c���|�\�]��7�����Q�(d�}Or��`ɖ��15���l��{eW���$ف�TJ����m'�7�s��!Y��I0��D@�b�� 裧�XN�����M�/�S��N?Yn���s�����S��\�����m�6���Z�Ƚ"M��s�=��w��k�6��U^V�⶗)���:0��K���9��R�5/w8t�Vp*��֬�RQ�2�*�x`�$��{G��{}�꟬��Tlw�`j��_��y�7}�u}��д�m�v<{��4ֻu	E�ݟ+��]��|��u�'N�|s���q�o���w	h���u�ƾn �7���j+sDW���@J\>�AFe�vŪ�ټ��=Fs��?�P�;G��1��5W����uI@M��J����=U'�5X�0ߤ:�2���q\_�Ѹ�3,z���f��+�ο'���U�\a��*�qM�0���]GF�@�~^�_C�-��TZ���%�4���s���`�Ӓ�)iחY^��)�_<
}�ݏٙE��LYpz��xb~a O�5�G˷i���/ٚ�z��`�Zd�7A�Nہ��F���/� ��AR>�}���x�?�
V��G^��YܳG|��E[F)=�0��m�	����[$��檞����z��4�+�5��٦���W�����G��!�|�����;��fzq{�:�>�3h�fO2pgT�L�qm��W�r��^<A&�%��1�5�85� O�?Zw�7
���L��-� N��=�@�,;|����$]SI�p�E��;�ݜ�
���Z�P�pX��O#_(��J�ŏ/�a�p�m�p_���������n;���[�{���U0UN��jq��ȢɁ�yC
A���e�B��S>�'����.x����:QO�j�!�� �,���<4��D����㠁����<N(�� �S�٫���94����m�ʩ��<+�'�fjR���^7��f�.g����:۾q}�ӊ!�Uru�����Ëp��ͱ��9������������j��ȓ�;њφ��j���(F�r�/륽w"7�cmL��uȬYQ�y'u:0^�K��PX�r$�Q�� 	�v[���U��^�a.���IN�P����-C[�6�˺Vhy�p��91Ku�#�,0�:a2le�٢A߹�!{{�`�8����DV�V����0�n����ZM|�L�h���.N�p��D�#�/��J��!�
�wsCє2e�7�p5�j��7j�*^ώ"��ȍ��d�rs6���Zgk)Mt��j��w�]�o�w��@�@�+��n���I(�|��~�{�a-��<8$�xݼ[򖺄�U�^��oG��v�j���l� n����e�� ���SnZkq��)@��<mע��B���`J�y�N����2�A0�hcvf���� u�`+��9o,����i��7��b�'T���_V!lJ�X}�T5�����Lm��X��3�;A�}�I?ޣ�p�o�p���x��e��n�P�ק�����圆�	��M{�o�x.�P�o���DU�2;__���iJ�lY��US�������Ŕ�2�4��{A��ȴ�zYY"q�u昝N���y�)c�?C�����^�`f�j�<�-\ؠ�e�_2�����FO��+����]��օf�������Tͪ�{�~�`��"#��1�r�5	x�p�ܯ�"�C������n� Ѳ9M�;�4�k�1ޥx�� ���U]�e?]�!�	��s���a`
Ǌ�3~���XǠ� ����R������'N ���?�/P2�͜WxZW��5�G�4i�^�����r����eb(1g(STr���5TA&���y>��h6�{�ov$�*E�֏U��%Ť�6���Ȏ�W��e1^fվ��>f��տO�'���ۄl��с<Ǵ��ܴz��!�?p���6�# 
B��C"�2`�3{U�Z�H�F}�ϯ�Z��G����t�rEFZ�W��c�>���W̡T�(����W���6-�l��`�jvHP�uEDMwB��J�j�.�{�l���~�Ǟl:Uk���xS�ć*\!ʨ��X!����˪�Y��Y�lI�uvh�`��~�22�c�%�E��L)@<��$���|ۥ��_+eg4���	��摹?y-'&���!�jQUe��J�f;P\]���yv�+Z�Zq;�\~��k�Zm!�1��Y�qkM��E���G�5
R���HG�ZE��.1�_�aL2U�˰����/.,b-�6�P蕭�-��t����0��m�f���$��%�S��}��}͠T��9
��4��T���o(B\�x�M�;0�&�A��%�e�o��2�D�sG���"v��]�P�/����&&���� ��_���xha�a���{fG��N�Q�۴;o�pդ���ت�j��~�0��Ͻ���b���<o��� "�g�W��/��#���� �=�$��Jf&�c'�:=�DP����ۚKAߣݖ}S���w#9'���̿���x��b��2��NR�ś���}4?��re�ÚF�k��Bɚ���%�6:۫W"Ij�܌�O��F(c��y���jޝ�'! $Hz�!r����[U���������MSa'��`j���Qf�3fb�9'�h{'�3��a�~��h�%v=z��w�T���7蘏9�q��-����
��y�uS�'~�T�~>���8􍨻�[�f�6���,vy�QK��8�%�f>���.�q�%b4f����"ε����������M@�s<�CW����k�O��xGc%���m�"���##��\&�Z����J�`�c�𒍿<�l���K���[�D|�2�`yk�6	��X����!����co�����VȎx�׆����&�1���y	e�.����H���� �;`d�0����^8�a�G}M�\�將����4(g|8�h�U����z��¦��僓�Md�f�m�D�ZŨe`����a��;a�m4䞡:�!����*$΋�2�g�F}�h��kZJ�
a�.T�L���iט�B[zJb��T5�JS*e�E� ��Ѣ�B=���W�[L������R�vB��k��'d�fB=��%�lnL�$��^���I5w(<�O���I۝�C������	�̽�3��f�"���/[h�p4�]Ol%���� �r�c���ё����'9�0��z����L�[+�D)���1"
0f&�� ��h]�6���3�L��m��*s�u�Е`y��{�x�U�od��mF�����S�B�ta> �/sI��M����2����{DZ3�]�{�S������-����.N��AP������y�S�asu �+)=�|�j({:H�q&{��<ʸje�>��0����,�=K��̑�D��,�|-s�<:zo��̡t
g���v��jE�����=��s��S=d"��*;p
H_�)y�Vʏ3S S Ǟ];$�
�s#" �O/�CW������Klw�uT�L��:)N�N�~��ת�J�AM�A��>��/Qi���Gbl2��^R�����uiV@��'�ϫK Y�jmݶ+����B$̘� ;C=�"��)�����m#������|�4u�����p@�%�Ѩ$��Ӕ����1������Dʓ���]�}x�bM��8a$ۿ>�c�_	��f��PCϋ�`��ޏjU�8�s�����梤랃l��w��"�}j�������]�=a�X��]�k0`��Tv~�L�X`:K��^��0��P{�r.�85��N�ߤ���5�<�5y�V�Q+����v�ח�ap*L`��qCS�(��`���(���RYP󮶇��4��_+*�g��_|z��N��������gp���ǃ��K�6���Fp���:��Xi|X��n��˴�}
���=VE�#;�03�s�i���e�����xIhY��IHRE;���"7�k v�[�o�R��������J�I`�O�* "����/7�L�OU�f�E�_��f�3}A\�X�CZ#Y��ys�����.��s�7c^o�#�A�r.缧����k�Ip��k�2Eu��<;'��Ò����M�畒��/F��.o1P�/����M4"�Qm�b����^o�ĺ�un3��2_n�$\70Z���C} iJ2�j�R�?P`�>�vLt�����j�aux�{\@���d�."�c�JƂa����Ճ��q'�/��"LB��9�ߞCYfS�V-<�]r���*�"I��Q���:�	�Y'����O ��` �7�ԣ�f�)ȗ(�_�E�Gyw�JjH�Mrw�$�"�/ßmd-C�F�	�J_�4�E^��I[�� 7��2�'��T�����2��F0���o��>s�Kƪ���+�TS/G]8��X�zW��n�k���#�(t��1��I�%20�'=g򾴞5�S�da $��n���B�B���+:����L��]��np��Ƃ��Q�`#�����Է�K����^i��%gH5QrV��b�wǷ�	(�q���Ŝ3�3��dv�!S;ԃ��%�P����g����8��@����̓���#;�D�`c�ɸ��r�<D�h��%���	�{(^>V3�Q��⬣�bw=fDSY��A�W��l)��E�#���&���q�Qew�{_�.����gYEs��������)���B��S�_Vq+��cҖ^[�N����܊̢�k���"8iaOZ6V����Ɋ�U�Oݜ�j$V��3㍥�4u�;�|"�n`�y.�۱��`�5�����}�~�4J蘛�9���n쨣���j{ټڨ�ɖt���ڇ�2��]{� �L[;�:ǝ#�uG�0�ѯ�M�_�'R���u������f��	D$�N0��T��:��%1_�����%�C]�K�{�3� �D�q �h�.�{���vZ�F�(e<�=9$@mh��q��q�I�蚪x5��C��B����0�E���3(�r0��u �m.34�K��	0>���`D0��/�f�b`ŹT���7n���У,`�-�	����E	��&��mh��L��� q�.r[3��GZA��=�Ʒ��XL"�"��z��x��y�س6�E��_��6{lsfx�����}Ǔ�_@穱��|�"��� ���:2�H~ɿ{����K�WE��ƋΤ�]�*7%��[{��:4�,Q�	����������e��� X�m�u%��Lݪ�[�eT�:�<����W��|��ϗ�.����5`A�i���׆�y�nt�LQk�9x��� �嵕2�0��t�鉅�qm�l^����ꮁ,Ǧ> �����4�<QL�zĻ��Jj�Y���e���cD�>�(���)���~#�iAtۢy���r�!���8�}ڡ�%�8b��7���Fo6�k� ���Q^�%�����~��^���J��,Ô���}�X��Cix�#;?7��,�m�=7Q��Ȓ��E�0V�aQ�<�\�qh�cs �U�!�k� ���I��f�m	gs��f�#k��O��rIm��\J�i�e��l�m�
H���E�7�|����B��i�ŉ��e�fo�X-���+nGn�.D4I()����&	׏�v`��)���4���'J2��_[f���i4�`�c��T���N��45 驙$cĝq� ±�O�|�R� x����V�����{x��O@��43l"�����=�Y��/�@����~�O!]��-�~I�XSh�P7�z�|@`��ʀ���F�Aս[���w����ƥ�F��h<�֫��^-��uJ��rA�@����Ut��4:�Ey���Y�Q����B9	S<uA?�aj��<��5-���O�	�Mx�C{C�Q|I�x�����A��� VE��[�#j�!%
R<C۽Z��l9U�L���]�tZ'X�6;oK�̮���V����^:Gvco��)�%Y��.!�Ql�ػvh&b��F�k�a=�?(m떣��w��g��粕���eQ&H���S-�#T^2AwT�-��4��:m�2�B�=+�<��nn�B5\�#I�ECI�
-����C���kg�=��=�4ǒ;a��߀R�1&ԛ�D�ع�ơ~/�2U�_�����
����>�3�����RJ�r=�E�MWj�y��a�t%���$.*���9���t��d�����������xk�� �*�U9��xmU����ǣ�����-�d�*�4WaF.��Ъ2�{�\d���ĭ���KW�
l��\��;H�6̙��k9�A�U�	D� 0 w��f�TJ�}������j�F<˷�3��N>
PC ���y7-���8��_�Bn���~�ŋ'����o���O�D?��q��l���U���+���ȡ�	�4 �?���V���C4���f��4o��ή[C�i��A
��X�v�����[ЖW�VS��P�3ڜ�6�;�V(Np�|�$E2"9^#Q>���Ɓ02GF�aGD�\E%m*�����X��9k�/qD�y��}e�3����|O�)�����-G>�)Ԯ�( o4�a�R�R��9�E��^�tU%�M��<��kY����ԋ<��3�oml\�fUy���i�u����2���ְ�h��.�?Ϝ����^%�U}Q��`���$�{�,-�{�y�j�&���˭%�"�	|ɯKRA�q��3�雤T�`"�m@:':g>�O=���/T��)����AN�#�N&�T�T��q{�;* i"0 T<��Ml��ӮL��%�)cP�T
_?6u�qS�K9����za&��-3�\�qO� ���!����o�uɷ��Q��KU$t�1M yxuǻ�_�a2�jY0�`���qxfPyY��s/�g�Ù8L1Q��荢uk�!f�AQ�k�)�4��7�� 1��*�t��nUa������خE#f`�<Y��)�������Tm� x��X<���X($�
k7����ez['�� X���,����;�`�3��)��������4aay}OM۾��u5��d�~mp���t�{�B1���M�Q
u1xS|m��,�2N������� k�5+T��e���e�5c��3;7�-��!p�d�ZF���El����p����'T|#;W幃��r��%%A�{#����Ζ�ff�}��]��k|��M4����]�����Q��O��[��ǘv4$+�0����{َ���q�'`����Ս��tCt����5憸�mJ+9�g���fy��D��Ty���U�v̍%Z���L�!D�u�H��'��]�����ßJ�i7��)���ā�!��������94}]X`�.�P:�:�R��P�Z_,B�ɡᅑP���~��5Nh�Z	VJ^s"��<#l�^���=Ň݈`�<��h�4ş�d��XOE�< ���E+�Z�6���e����*�H�|椇u4㘛j�d�-�}o���@hF���)�HpU���H���t�'�nInI��\r_��K9�]�ni��r�'6_�la�C5��i0�� ��\�^�y�$wUL��:a��Ԧ�u
�#������_�_�F���i�KQW�X��y~�dRI#�ͩ�Z��mw��<�ZaL�M�Y�d�M�&���R�q�ψҷ�2�a�#d�1P�.Q��ޞM�[�zqۼ14ld�����un�g��(}O3��B?��z���"�=�am#�)2��������z�[M<~Ccu�2�$�V�r�t�-퉙�=r�q���\�Te�g,��hE����+�ua��W����cDi�lDk���c��6�G,��b��k�F�x�2m1 �F���fxpG����/���*�W�l@�A@
c�4�OR���}Է�_�*��왍��H4u�D��d���IO����(v�w�#���L�<���� �1[�2ъ�uo�V��1\	�Hd5�C+ҟ@k"�DV8yyd��j�WMU��"2�������N��hK� �BS0t��ຊ��qQx�R.���]��þd��KR0�g\��s��ک�`���8+��(��Cl��G�m�#m3��ȉx�As�s��_q	�[�9V^����� ܗ�-����� �kM�8\�������������`�
���xK�����i�޲�l�w�� �,?��֟"�Hz+�;W��ClΩ��3����wi�I�q?U�nxa4~�v��g��iMЎ;�'�3��?�(D-f$%��3nusnb#b����@����Q�����]�	1���C>^��v_V^#�O����pO��A�"�	�T���"��Y�P�����~a݅T���Cxa�q9�U��	w���/~%��QOJ#��]q7Z�a�M2��B~۶!Wa�s�6�IRY�4����9�F���.���pu��c]8?��hރ��E�!@��1��M �ǲK�����v�9�h�!�����D����V(T��*n"|٫�
�I7��'�5�V��l�%�/V>[�v�}Ij����Z�0�(o���{��*#n�3��R��-�UR)�g�9�]9��4[�D�[?o��FK�������O����i������oD�)��A���:ڑmӖMa����A)�(��r��iHh5Q`��D���*�ک��j�G��F�W�#z����Y|y���,��ñ�n���5T�Y�j�6O�ޙL\�n���I͉��ݼ$s:�ڵ�RJ�����������#�����l[�o�k����^���s��-�
=�2a�T��qi:�����rS"1�p�FC��T�U/�:u�z��$���huϗ~ �DG�t�>�Ì�(�#{�VǷd�V�H] ���Q&��VGF��n�B�;q@�B�t������"�P���aT`C�-�����Hq\zR�L����ԅ�O*2\}m3�� ���P�u��F�Ļ� ���1;�r��V����d�Ma틸A\).�bE��J�O�u:�b==�R����~y)CnD<�a�ӳ�����=�;���K��i���2���2vg�&k��8��X"�,N0���܋��R��� ��B$R�t�x��{P^�췗�9����T{��	���Ù�0O��!��e^��tӝ�e��Cы��a�*�ۛj`��<c�\�W-��
+`�zݬ=��������h f�ggT�0�Z�H����z%(Y���ѷ[�w�M��l�T+��%9ƊAB�K;�ܝ4k�| ��c݃�d(TRs� O���4k������3������ �ܪ뽧"��
��h��k�����S�A��~u�A��=Las{S�(�X[H�N;Y�"��t>�gKw�靮,zY���G/gTTVY����x�EK#�X��s��^5)��jmM���7M�7##��S�r���F�$$��n[�wp�<��M�Qyv�ء�Ȭ�V�U���p@Fd���~D�/�.FvHy��_ ͜�?�	�� `�0E>䴥��@n�=�����p��0�B��~՝�v�@��B =�yb�߫G�r{������'�勆�#�m,~A�E-9ꢍ�P���{�-��ⰺ��Z���E�PBt0���e����=ʰ�����A�N����N�T	� �o��4�49"����Uy��m�qB☀�tI�$��Y�St��]B>E�����GR)A���j��Z/�J�P^�KP���e����]l;����ӫ_8�iѼ���<ӊ�b��<%Y1�DN�{�K�?y�	�����[�Ó�Κ���'Db���yˍ#���JuA�ν�.ȅ��?�M��r}�w��ǀ{�Uw�Z��*���7�+䙌;�A�����hJ�z���l�p�]�$4�pM�sW\���2�YnB���1�v�(��¤��Έ%��Nhڡ�������+�^f�w;����ɫ]�eV�X��z��B���6���t�E��v��DG�M������D�Ƅك�n_�ĒL/u�U;�φ� CM74���^�^cҖ�_�,2�CY�/(���x��@bR�[]s�P�]�y�q�]���7r��aB���:S�����L��&�R��Mj��c�8d�U��j
YsRp T�b	��L\@�,��M��3qcLf�(�N��}���*�T��MT�j$n����cIs_��hb��k��&��^Q��L��'�Z�AA�k�K��xEu��vsӜ�!S9M� YYg��X. �q�uf���U�Z珷�%h@9��*T���_���Q��gyڱ�ޙwG�7�\�5'a1������gw�������,u%L�TB��6�Oq�778�T3ڽ]�����u2��i�V�Y�ɽ˙��<����(�O�S�G`Y��Ʉ�]���A�|�A������x��ɒ�'=E�<���M[��^�6�|��v
����>G�#?r5��\S"b {b����K��ȘK�ߤ*�>'_=0�G mib��l��?��w�e�'a�g��fwr��f8��\2{ TW��i�+���_ޝd�k�䡽ٔ��L�����{�3sߐ��4��E�%O~��_�z��]gȠ��
�_�z��%�m�����c��0<Im��0�Qj��-7e�?��S1)i�u e&q�g�~���:��2o D���[afvÓKp#h�A9Ȋ��lB�)�2�v�SkXl���HX �E���Le�"��E�;����@�*Kp��I�ǈژq�E�P|l�e;=�C��s�LL\�鳢���jx:ZD�7���j+�b�KB�.����A1�ī0���D�\��l�t��Krw�ČO@�c?0)|��G�
�B� �gU�y �G�X� ̬�˗��"��n2Nd����~}�c�O�J<��)��Fu&t�	��Ƒ��]�FT�!�ȼ�U�C�n�;	����EU�r���w�0Ѽ��z2:��INӾx��Z5p�'�X�(��V�����.�ŧ���g�:fܾ���>qL|�)Q���X���^����ԜP�(dp|S����ٙ��">��E0#���趸�}�1c�Y%c^}���A�^>�l&�u��|̀�i^rN�؉��͍Y6�0N"��$^�cz�r8�n�������A��{B��	.*)��CZ�p�b�A���������.�|	��dB~ɟ��u�:�c]���l�~��Ϳ��pv�5�8ِ���|;��]��s-%���9ڎA���?�^��L��!�)�5h��D1���e�Y]!�d��yf�e,���/�j��d��$��d���
���46�_�ݲ��P��a ��⮄P���75�Lc�>�4mг�[JH�t�> s`Γ�~�T��)x�b��i+�����8��	�<ؽ����_�[3�0�/��S�\4����$=ӽ@�=��� �0�/�p�8u�W~k��Ng�ۨ(�Fnq^܇��Wx��mJj�e���G�HMl�
�y�g��0��7
���S���2��ވ�Y,����b��_�?�T(,�	tnF'1l���x�)�D�J��I^@��|���}s�^�$�=d�7X��KG<�N2�^�#�֐����1�W��c�Xn�~_`�apٰ�l������%�N�j�moz��t�ײ�>�3Eǈ����l��.$�Bk>M��������,�t�����-7&\�N��E�4���H�:.K��n�E.7��<c�3`)��".{�9�U*���Q�A��ک�Ӎ�ÿ���d:T#
��VO������WW�I�������{�-��h8rО�����i?�}����΢�on�'0\���7R���5J�3ǥx7Q=-�C�x���	�6+O�yuxp+z�����Zur<�{�e���dt�pK�D��VI�\�E+�B7KgE������'�X�a�3���d͠�|�a���JlQ��K;P'D���fae�XG�8�*�d��R���`ur�B��^���ԧ1r>����*K̻[|i��$#ב�u��v�h�KL�\!�?K;��ܪ̭!,L��0�P2����M��	���<W�]P�7]�=Dz�u|�E3G��@���DO?�~7�k k�g1`B�S�ε��}����"x���a>FB�#xa����$�D�q�+T��V���,2b�r��O�^ޭC��a/�Vfq(˄�Oo)!n�D2�Ւ��z��t:�XW��%�3�RGs��zv�^��:����"Y��̸��ٶi�1ѱ����B����|1�h�e�>O����ݮ�A�ζ/�T����}\1��Z�.d~3c��#=V�T�z}��q�I�˜�Y��>߼�C�?�.bw�9Y�w߰����!�5��){�ɱ�dï����|�TV0�wQ����3	�\���h-`��������~�R�i_��v:�4QBg���auV�,/y�E��8�=��G�\�E"��8�=�5�ӈd�$E\)|�{Y�b���|��Q΃���(�Յʡ����c'υ#AD���9�u�f����tV�&_S�؆P�FB��"��?.�r��Jz$�jZ�Ѿ��DEj�s��}�Ă���K�����1�y����K^����yU��,�f�eN@�TD�v=i������!�.�p
�,s~x�Lw��& Y�ʩ��k��C��T@�����z�*[m�t��&@�pXp�o� ;�ݢ^��8��[� �=Y���8e�r�G�x��8�=�N��e�����O��׏'�K�]5�ǰ����%� ���)A�x�W�VＧ��H�a�j�w�+0���� τ[U��ܺ��M��D<�)���!�bȞ��zt��K��[D46ÔKow�2X`�4�)��9g2�P���p'�z`�"�	���1��`��D��������+Q�2�UG{	s̐������Yy �T��� ��$W�XT
F��Y�]N�J�_*������a����vM�P��""F��2��?�+o	�.ↈ���_,���<*�6��2p[���/�(#`�bk��q̙����0}<-:Y�q�2f�zrF�@j�������6�2mݯ��
�˔�<�@��D��I����+]N�Q�˭ŉ����i����G�"yLKnt���� "���KP��5a��""~�T}��:_2V��ܢ�+7(�C��'9��ӟ,��Mog;:O���E:�������^0<�Dt@t.,k�T�u����� �ջ�11`��tk�>�/M\E��<`�Z8+���%��nß�K���ե�\����g�1m�2M>��2��">�p2:hD��6a���x�DK�3���9��莦{�u�7%a���=YGQ_�iťK!z�CXX����أX��"/I����2��KF���pu'��(�K�u
���T{���u7��j�t�Y�G��/��B��JN&r���l�,�ڎ7��R�!Y��L�<*�FH�(�;��1���E�\��'��"�{��� ?�.���Am�+����#{ �~}7�q//�|��#6!1	��c�� ���;��"�x���t�q=ṉ]�Z �^�&��4�3�$���a��po��u�����B�.�e�.x+�,���|u��1�.p�d�m��«�jd��Qϳ30��vhL��ӓE�#"r�X�+��	 ��Z��#�͹�Z֬n��WeU���'R�I���ߢPF}�CG���ƚ�؊<�=�<e�����8D<J��LL٠���T���c\�ދ�.Gm��[�+,{���׿�FOl�r�>�!2��#�m�X;��A��d/���Ȯ��|`�ٙ>ξ�Y���K����XK�x(;���Ї���D�V�������d�Em�^dg'HJ���D,��/P�Um��Z�WD�s~���������Sl��3� �Rt�XFn{-���d@w���\J�������}��='�yپ��[�tgF��!�G��yl��"<���2c��Z��ħ������}gh�"5X��5m��d�H_K姼��y��$��U>_=�Q�qJi���������E���44��d��V��ih��t�a��_�w��W%�uJ ����~f=o#����XL/����\���6��!P�F�$wv��ǔ�"_�
y�΍_�-�R�z�K��p�3a(�'��ZMݎf�ZY[��c��>�����~�ܐS�i}DU�y`��?�!!��p-�'�Ȩ��= �M)]Z+cf�EĺoF��A��c`�������*�B*���7H_:�#�����L�Wc��M�0@�P�]\�K5κ��{�9�K×��!q��^M �n0����ʞ�X��:�P�<�z'�+������P���?�o�Hگ��G�����@�05t��̙�_���A�Åy�-�\�(�DM���� �%q��c��b\�9�_��:����X�o�|��%��#v�d��_���nR�S�Ъ��[��t���ƈ2�>樼{`as�1מ�4������$g޵��8-��٤<��Ϩ�?��㺄E]d� !�EI�"��v�.��Y����~�fPC�x����1fIڱ���'�wo����$h�w#�K��` #�6���[s�:�ƦK�Z0~U\C:;����|6�,�Γh� ��Z��'	\r��y�D��*���8D�����A��wɵc��?�Z�/`r#�G[m5K���|�/7�j�yR����
���~�j!�ݠ��2� +�G�b�s"��C���c��i�D�%����Z�$��pf��ְLA�z�]Y�\��ǆ5A)��aZM��:@������[eg;��� }�z8>j,̇@z�M� 49e)O����H���Y>p�\�b��H�-��S���3c	X�a%� %����Ӭ�! �P�^1�}<��	���&<k2����s �h�O5��$s�-�R�\#[C׶-ĮD`�&X 
u�S� �5��Ȼ*13�#�/���� &KY��:Ȟ_�,�6��Q��)?X'*��-I�U�SW���pbژ��-Ճ���j�.������?[�R����+��p�ȴ����2�=T���������>�a�����UArU�JY��~'N���0�I��%���Wۮ�|L[G�غu^�,)xq�Wq�L�T����t��i*e��w<U!�D���K}T�ڞ]j�_zQhq�)'��A]w���ଏC�Rlb�'��3@���n��7�6��?��};f�J3-����Y��3�G��@z�sۤ$���O��b����������ÕY��ơhW���o�Z��-� gpk�sn5!�����ζ]��,M8\G	��7��6�۶�^��	���^G0�����ɇ"�f�&�����?����)������n�6_I��^���UD�Y�DY�"z��Ob �0ߡ3:(��! ��Q��x�nK�f�{��4�$����C�mjz_A#2����m��#f����\�؃��aQ�}LʲM�b�����j?�3����&�Ի���� J�����@4�(m���],�2�4�Ԑ�;��C�y�̧��^�s`��]��[%9uqz�L��Ⱥ�	w ��:�k@���u��B֥y�>�s��D���ӎ��=4Q{�"��������1։pF�g�Q��: �ֺ��@�5��x�&�,J�T\9�0ݸ��\��4݁1�^�up��.R�� D΢��yM����I(�^�t
PZ�ej
�.�;��D�/zV^% �=��=��1�;aM6�Cz���S���|��A��5"h�1л�]S� �0`9�
]�i>�f/&71�3�����n�����]E��	�U�Q��m����:��_���c�h�̘����Y�/�p CP�Og#Y�?aQ.}��D~�!�/��"�� k���� ҔC��g�U��L+�n<���D��c�|��� /x�_��aИ�r��^������e��H���ĳsP<�H;��bk)G�<�$�W|/�N�`/�o�DH���Q7oC�p��Wq|�o�f#$>�`����p:U�bH�@���\m��'�݂Ă��`=Ue! },��v��,��:�ǅ$vkX1�h��%p�F��Y��)�Uh��$�jJa�~�h����lq�Dm��f"LP��0��t�/�@�%���X��4��uw�F��\���4�1�4U*���m��e�$�	Σ�H �����a�H_?q=�]Np�Ϥ.�J֐ïm�<�EmTh��	R_��h�|����p��NJ��n��Hcb5�C�g+CY�����!��,CZ�񹝴b�gU�<����y�r-��i�����&=�3�<=�)�'�$�4�hW�W�[�n7N���,b!����}��_��9
92�_N"��y������"ҡ����V��z��v���O5��o�����W���/xX�\��8����$�s�m��㴨��6g�;z6h,l��::�����N������:JY]����tuY�<VWl��/-��k��ю6ͼI�%uZ�pPZ!{4�����WD����]|��F�s�wstc��B|_BT�ǔ:�-��K.��Q�̈\��=K�q�D�"��g�\.�D��ý/���Q/�5�x��Q��X���I�	}�����w�B����^������s����/w݃^�Y�m����%|�xo����* !ز�MӼ�. g�W�<զ��%.K�#��wG�i<?Ì���7	�3��L���q��!�z��������� 8qu	C��_��˯����~X猘����u�fq|�o �o_��6Y���΅�n����xq�P��W�u�>832:��OM��at@3{L_p��On^�����`�
#�X,�"7���M�3����b�}l�퟉F��J�ȑ/D\fZ-��T>!��ð���Ѯ��_~i,���{3�"���8qT�@ʝ�+9�����Ԗd��iJe��o���h�����c:���V����\��ݔ������ϴ۱Yh�N���bV=�/�H@r-a��I	wW
(����$���=��A�eK[���S�4b��?�m�)��b>D��O̮ϲ��'r>F�9�zkr��&���U%����%�*06������ ��ײ,��ފ�1"���g�<��qU�� ���+��R�T��pY�`���|Fǚެcj������v�k�\�H������?S�����w��e)8#��	հ��iy%7� �H��H�o4\�x���^�$@gnr�;����=�<��ޗ�{d'G�/�D�}��h�AZ
�[{��;��8��|!�pg �P�]E{��6�n�e�U���^AY���-���:uY��BbZ�U^�+a�\�KaT�p��=����v��O	`b�XsA$_��5"ɕ҄1o F�`��ܳC�:гT<��>��+�� � �� 1���t-��G�z+���}7dx�)��}������Ԧ�[?�d�_r{m�aM^蛆��}�Pէ
�$�v��.$�X����?�(u�t����Ms��}�o��.q����&�O4;ݥ��?N�	��{��BM�����T���0P���^1�=N�̓�mD�����&<���	XH��� CkU���Ug���b�N^0& 
�p�٤�[���@E�JO
�X
w�.}�gIU��Ī���	�:��ъGx\-�Ə��Ѻ�P_���m�i�I٨/���:9��
�;P��pǥ���ߛ.��􆩢Gǈ$��a���A�<WĹ[���d|���fv\T�p��%��`�Ӈ�hFT�D*j�Ek�f�M�HlS��:l1�.Q	y�/���Olְ�Vs��<���!j#sΘ�~�z]2ލ��bE�Ͼ��d3\�g&��%	q�����;�${Ȭ-�8�o���6Ϧ�)���z]�r���I|}`��Yh��?��z������s������M�BBf�o5�K�E=��/_]�+�5�Rm���'��r�p�N�0��f��5vEbs����8D�>iF/�A��M���/�-� 	�K��*O�A����!"���o��9�H���5s��c�[G�P��ޒ��?�~?�j����{�Ӑ@BVͲ��ڪ��n��Iw#~2n( v;B/��T5xc�<Ӎ~R����p<�D�#��z�Õ����Ę5V,p�3�� ��������f�#0�WwȥG7�wD�t��(�]E�j���<�=��m�>̯iA��;8�Sk�Ֆ`��_��)l���)�TOưC�֬���O��x��IG���� (��h[��l����Z)�Ck?����0��'��}V�lD,/�r!a��f�]�A/��Rf��f5����eT����,�{��o
_Қ�z��3-�~��H��������9��jg�]:�6��̅�U�?�A���jU�䞄�P�4}�x�ŋ�u�H�9F} .]6�
�e�վ�x�d�I�A=�϶���qv�)�(�L-(����RQ?�_�$8/̧��q��h�Y�ؽ��o_�(Rjo`лv^b��*�r��m0�q����eR�SZm&c�0��$,� Dħ�����n7p~�>*�	�d��kMt\HR,���H�� ��_��q�a�)Om2hNhڞ���.�H���{s�j/�{�V; �E�{���E[��O��V�ފ��`���]I;��@���Ĉ~���l�����e��A-١G�g�h��w��R���@1�,>�!��Ca��9�S��8I$Y�M��C�	��p '���dZ������a�J�����2��n>!�[��vSWF�l�W	 �!4�?�߳��������-	�oCB��6���P���n�p���Yнx��N�t��A'��)��Z_Q��,���j? �Q`��%de6��M@y�a��Ar�,�&�IE�v�љ����~.�x�?�����S����џ�������z)�M�-T6�@���R�hL?�S�����	_y˚����.�����ݪ��7���>;�Ơ����i@��٠� 	+Ok���q�Gs�F���Q
]� ��3�AXG�zy�%gyp/�B���AZӲESl�E«��y�vM��6$m����=�h񽝭#IYU��1n��d�Jn$��ܧ���#16~��޷v��v,�H[�7��ipt ����bqG�m�`Bh�wjj�[w��k��L0�B"�y3r�
;�
�go��J |���%}\�Ϙ&6�1r�d��>;�X�eե�B1�Z۠�^��df�T@Ic>�2�s@r�e��EKߴ�|�s�OG9s/I(q��K񞹥��=PN13<����=ER��u�57u^˓��e��"�'���.��흣��J��x\�d)W����+�<�k��e�yD�i�c�J��WE�M���_4!�����
�k���H7��	_���V�b"g1T�X�EN`�[�Ӏy�@�I"�fK��djk}td�?L���jN5�1�����Y2�c�cb,,��5Oll�����W�!�@J�Chd��|�lA��e�)ME^�]I�0�ĎDV��W��@�eGY�<��Z�?�_�%	��_�_���Q�ª>�ƨZH?���ęU� ��W,rD~ �G�T��{��/'����f��<)��m�r�Ѻl�U>�7�vH>)�(h\�y��\jb8w{���O4'{��>|�-9ע�
P�R�@@�le �9q�2��� ��4��3>@�X����oRMe������inxYz�_��˟<��%O���װ��߬M��A^�-P4c{F!��@T�dk�����!ѯ����T���WP(U#��MxK���N�d�|Y�?��y/���U7�A���6�V2�WH%�ĳ[&�3�w'��d��K� &1
�,1��[�u������^/�YZufg$D��	�6i��o��?�7��Jo$����47�����==1�)$�0�}m���d��2�m[�d/����
��W���yx�A�L��t�{��'�S�a����1�F2��br��ŮU��"���,`zB�mB�����͕�#���Cp�_-"�i'I����{[2�
'�GP�����q`��]�ѭ��-e��3:p]�b}���G��!�t�ל�#]W�n�u�"^��R�K������}�d4q:>��E}��Ow��A�)7�m�yٌS���ݍ�^���f:k�sXӄ+i��	�$F�2Kk���!C�]��R3/)R���j��jT�@�9!@,{6���3ҝ�C@�Tr��Ǖ;��A�1Љ��/�Sf�����W�����R�t�"��t;BE�E=��*��a��"F�є�gTan���^=��N�< �#���J�6$�0A�!.�kP����A���l�Y!�b{��K��dA��$����4_�q�î�5���O�C���z�eW]Ls�U��x�"�lB�&r.ѷGą�`�**���*�A�6�B��j�Qh�X:Z&˗TyhD�@��@+ۨ�o?�c@��wS�]�#3��u50����x7�	�<��Q����^y��L�iQΛc�Y���Ď�ŔZ�͚d7U4Jƭ��bcު���Yx�%��ƛ ${U����:���+�k䚡�5�<��K�7�̸�w&�ޟAiNI��nK�r|����S�-�K΋�pmn%��a�*0{I]�z��er�
w�!�E�Ha��i���jN�����_�.�Pj���m֒�:c����G����k`]{DY�����o&���gv?��A�?��w���F�P�錘	�I��'���cu�_\a]��N�
�k��`�TX�X��s�?!�y�����Xn򗄄�»YwS2��|1ge�{��0��Bݵp���������XM��Îv�x�iDE�5�f������Է�D��K23ݹ�K9*�w4`����Q]f�Z�Π?T9ѣ>�]c<W [g�@���D�0�ݫ(*Z��f��)^��QhG���yR�RK�٨�D~:J�!�CF]�$О���Z�A�Ӣ��}B��Yն!Fn/�)� k��1�C�-�Y�te2Bk��J�)�G,_Po�"NzE�vY��J4\t��2��2�a�(������a�<&�7���g[S���<wAR>=l
�^ػc��f�g��)�m�n�xS�`�CM� ����$��ة��e%�>�.�#��v"ʳ��'b���6l���sX���{��J�����m��$,�1��aQ�D^}{�J6���V>�k8E��'�]B/W6���`���uqfn�g�����$�71B����o�\�d�ϊ�k҈녁#����&K�ϴ{�W��&`�< >��AZ�->���^4�yP��'���S~ȳ8�=ʵ,�8U�"tP�
cCS#�Ѣ�?�-!��}�ޠi ����QN_�{��7��#Q�vpV}�;�a��1�5�t �����J'�U�V#��I�s!���>��5�s]
�=���G���+ww��˹��9�
����T�Y��u�s)���1�C��|�,p�'6��q��e�~�4�kb��G���p�wTR��R!���>�A.U>�Aǋ��ѕQ��R�}g���H4�Φ����(x���Xw]J�D|mCZ}����:�2vۇ��i�B!͠I���f7S�$�jw� &�����3-��E2�aߑі�� V��{�kG��_��`.���\�,�������J�7��z}��zN���?�p)�pt�k��m��*��c:������
�]bןJiؤj(4	�C����ю6���D�2@^T0+L[t5{�ք%�v�$����I�U5��.�PA����5X"���7 �h��T�>�iM��)��F&Ul�ջ%,�d<G b��1�d"�^�,B	(�á��\H������Ts�Æ�"���\ܝ�ټ�����k~����)��"#�1~�g\�E�Gޱ�i���#'���y�@�Pi��u
}Zx��(��|A@yy����(��f{ �3Y��[���ƽ��?����4|\r9��l $���Uz&=
󝽫�E�L+{͇�����lO��Ծ���[�������E�c�]a#W����M����*7���0��b�.A�Ts���6.?�
�>�u���N��4��Z*V ����w�_� P��x"��HH) LxO;H	.�qZ��߂޴:��^a�=�{�`��k��K��KzA���Bs]a@�_H�t�|/�Fr��ګ���UEA���i�.��߸�M�����$����+Qr�E�]�u)���<:���!�N��0YUU��Y:lg{��u(�'���mAm��U�M��o�h��Fi@��' ��l d ~��s'�x=��"�D�1&�Ӿ�9='�����h� `[tb�bn��zc�IM�� �%Ch����1�f�(�Է0Jps������3�׵��w��~��{��ph���
��,h�o
���7���%��d����&m8�q3z�\!�t�~KPY�
���J�n�����Pj[V���a�$Y{�q;]Wa�7�����I���*���\�}�-;ǇqDju�7��t!�=�Qn�nh=�n�����-���� %�-�)I=��Ze5��Z�՟t����S�X�\�IK���һ�Ǚ|����૖/��*���:L�&e� �aZ	�s� y+�V��2��M����&w���X.ԕl�O����!�h��:�'�H�ah�w\����K�c����#c���?�ג������M����`�X��]� ӎ�&�D�'�nxq���|������|)S�x͇��QȧQ�����Eh�>P΂�D�}z�v����$��jj��� ��_���$E?&����Yg����
x ~�jy�5^� M�^�nuS��=�m?#�m@�h8���yl)�-3��ݵ
:��`d�i�r�����*N�д�%`�\�T�N����"��a�ߤ�������k���#)U�8�R�qf��*pb�B�Z󦜔@�"�9.�Us�T��-���88d�m?�ei#���`�E�>�w
d�CQ�V������K�S��T��lϿs&�z/ ����n!�6*�.C��>��+��l���<��/z���-���S������N��[�/�0E $���=>�y�a_3dT 0ҙ�[מF����뷵@����V��=�lj&��hĨ����5E������<Ѝ�?�}gZoO���ي�\^�X�;ߔ< ���Һ̱L�J�t�`)X�Pۛ�9��٤ �0I�I�$�C�-�i~>�/ieI"�_�I�����wJ���$'��#�ȡ`�p2���,a�Lg;����n^�Ǣq��+0:(��ߋԘ�L�_���L����l ���BSԕȿk�5/���6F;��Cxk�Y�y�:��2Wr�N�gG�6'~�L�����D�:�41 M��2�d��t�J=<�`GQ�/��1��G��HjE�z������d��v�2�"��F��2�����g�ait�I��,8?P����f
��ű'b-��*2���
+界7T)�����7��0.�\fq�9?���Y�v ����_$�;qo$�Uc�W�V2�Z���A�;����� ���kّ�lVV�cp5�� =���AW�E5�5񑹩C>^�{Q��!TK�-~�Cn�!I
7�9TS�֐*�u�ПD���Ȏ�o��u��p
�V1�s!"�J[mh5����ut�|&�U��u�T�4�H/���C�%]�n~
��V�&F�t��g�%Ě��Z=����E
$�wun�fG�d��A�j?%�Oa����)CM���h����S'q��˧q��?������@��)9�7ٗ}!�%���k�����%[.��e���g=�_/�k�tiw�x�r��蘁���U�P�`�՚�;B͏��n���-�!;�MD�@C{��r,����;O�r~�{����m^1����WDj6��b��Ȕ����"@�	3�T�~vr�p�M�:�>J��6�y/� �a9HN��u��M��'r�E}��Zu@G�~�̻�l�L8�����|�ȉ�\a�a��@ϯ�{(_�J2o��Է'�UW�O��20�2u�Ѽ����ß��bQf~~�:#���*�ӂw�?XX(��]���)�)ŵ�!�¯K�_���+3���ij����.��Q�*�z�8��{8N�F<l�t���Ɓe�|%�.z�����|��?��M-�!K�2���ק|��1�X:֍kjB(EI�_��qy{�}�������!���'��IH8�<��
߮^�wK��#���R��4��hD�
�G��TN`��W�ګQ�_,���HMO�ac�9�r�M�,��R/��R�FMN��m�$,��Ɩ��G���U���������HH��8�:5��|u�J JI�$&�bH>�r[�n �̮��:�i�e����l��^��sa�,���ӦL�Y�$�km��)j����%�6�*mv�T��̀!�3Iw��"������m��/�r�m�(��n?l8����|�����ۋ[p���~��h�Z�ɖ���9u�����r����.��}�\�[E�S��B��?$m�8E���������{9� {�FѷK��ŒFQB�)K� �A��'�5�U:���-�z����F�Η�2ⷩ�7�&R�Y�t�@���Iw�t"_\R�.-�HW�<�V�M[��A�l�X� ?��)�~�b����Ѫק�̲lm��̤��s�t��\vnv���M��R_��������-��V�܎d�s�O���*�����}J�.+���n�ru��|��y���J�L� cΕ��1����}�.SE��J��\ne����wG�r��373��.́w	3��ŀ#M�����1y���A7K�{���v����Ju]���ʸf��څڣY����]srOp�Um�z�G�����5ESQC�擳u1HǚUi�\cQ:�}��/#D~�E�_x �C���9�6Rq�9���;	e�Ly���^_{�j���<�������A��4���+��_{�.���]'���.�S���ϯo�� ����X}*�{\Nnͮ��?���K��RI0(��]_ዴ~�h�����xg˱���}�1�79C&�P4��a�rG�Ŭ-�X`��"�'9c��hjF�9IGK��T���w��������������C�9
��ù�B:7/0:R3��^�p¬9�AKN�!���׼�T����t�d�.��*�`����V�� d���W�U�`��Z����mV�'c>��#(�ԫ�qq_׵�%v(�S���q�o�+�Q���ަ��U錊-4Օ��w~_������G��[���`\��2���GZ��s�Ϳ`8�h]���Cʓ�{�3��x���с�8J��W��U�HQ򽺤&X��!�lx+�.lZׁӋ�~!��FtM��qhy����S�A�0�l^.<yK��GJ��,[]/���S���>z�#z|�w3���Hb�1�e�kT��!+c8����dj����7*||oz�ک��g&�(�w)��a����EvN��ruF��@I�7eP�5W�or4Uv <�s_.�m�R�7���P�9�e׍n�4%�U����H�u��O2��VM]|�M�թ1o��w8�
u0IU�/��� <���I��l��}����J[*��:xQ]���0�
�����(�$�#	�tJ��䤉�vJypϡ��߻֐3�����& �A���Д���\�tC��/}8�Ǎ<'�k3�?�#�.�����X��юS�`׽�	�R�ʫC�>+*4�8���<kb�����O�RQ�
�6Z��
���LA~FJzQ�t�7Ų=��ů�,�|"��R4�:�Y����Y��ޜ^r�L�����j\��u�z�3R�����y뚆��I��m�[l^���j��{��TUQ�BH��G�!_���3М�&�|"�2��^��(�?
��8X��PT~������ѽ�N�4!c��8�*s�x	��;�L >��-h.4��K�[����o���=j>�5�/YU�e��$w�U�S�ߺӫ�gT_YcCk� '9���`)�1|� �`)�i��x���uX��A�!�,������.�)*9D�#TW���B���-[�J1]B����F����==�ޭ,�5\Y�hA�a����C��ϙW�4��Kߕ�/�Z8#9=7{97����,���Y��<�fQOk�D� ��r�i}]��&�ny��?߿FL��"mO(x�kq�j��Wl�2��4�L�JV�o�b<${k���ƦJ��-�ݢ2�oy���6%unT��}GhYb��e4��g-�G'�������Z���L.L�B$<lT����Ex�*�,�GV=���u�^I�)[�xV9ݰ��ND���l��-�>w��V�Kh��?<���6慟d74��V$�L�A�d��YK<��� �$+�����~F����a�`�6�kƘA D�<�([��*���^Q�xF"+0�v��d4�юژ�#�2���u���aDd��-&�°$�0s��]�A�߈��e��"����WO�eI�@Rv��ui�a�%��R1��1��蔢����]wm�ޱ�hZ-q���ן{0h�懽�4C�Q��]��'S��� \5�/ƞ��a���U��o�^S�z��-AJ���Y!ۤi��t�SI����#�!�IfA�B���!�� �Aҡ(�l|�I*Z���]e����3'J�,����9��O2bB�z�qF>EL)Q�y�R��c\>p#�0����Q E�΅R4(��s���5n:)y�0�g�m��|��1��rɟo-L=���)����x��ZΛ�u�è�-�C����~��'���}��ʀ������~H?�����/$��gm��ww+m����;.�vI�N��!*^�0��~��ݝ�߈���%>�΋l�o�;S�/t�����&���};ҙÉL�.�ܖ���Ti:V��_0�{r�Ґ�������i�U��/i��9��>�@��	������3>m�>s���_��}�)�<+�D�m�ڛ���)�w.}ȀpF>}Vθ����H�h��Ͼ�
��])D�n=��ډ�Ӭ��Ը�Ƨ�@v�)�GJF|��J�&�)G"�����^��Np|"B�\��f�'��Q}�x��Gu1��q�/���Q^���8�THp�"ja~�NLt�.���V����i��t	���d���0�&A�-���ɪ�����|�-����sm�IE�-���6�����6q������v ��_R����3�su��	�f�D�hA�h1JA${��e�gx�꺨���1�����w��cd$`�x&k[[���CL�Vߝ��zK0����9�\ĸec�Ơ��t�)�P�n� �/g�Ɉ���	[{֑�2u�ެ�.G9�T�iȥ!/�/
��N�݈đ|�w#}c���>��w(�r����)���}���1�SUY�B�@Z?^9���JW�Ұ�ߕ�����R�5l�9�Z��	�W2�d՝�����/��F�N���,3$���	3k�ͧ��?8%0���iM�i0]�`*��=����rG��%cQ�L^���R2C�:���z�	�B�.����2���鎰}&�I���YN��O44�_�:�

V�E��Ҥbf+����ްè�|4'�mAG��٣�J�Hq�|��`ѕR��4B�oʣ�iB:�$6�Ȏ�ƏnK�Zj)��:<��{ �v⮄���B{Č%ɡR�q �ߑꚝ�T,8�9�8�7K��s"t��"LP��_\�<gA{N�����#��%-6|&�~�F�OM��8k� ����I?�U} }����*tDBT��!����ɣ�|�A�W�}I��.�ٜmo�aXd��YH�j�*��}x��B�'�Y`!�{atO��w&�b���gV�;
ֶ*蝐�Y~/&LD�D8�&4��;� �=��;h#ע�x8�3��8*�
c�Z�F�Kx@��A&��el)%��MCX!�.��4��
�"���d���*����Tn5O]�v����������A�d�b���~�{���_PC�'�7hawfP#�`g�}&ge��)BN�ˤ=��������'N�6�J�tB����>��oc�2UjW�<�U�t-�9ceuSK{�O�����r���j3.�t��?�/-l�5i���ǝk�C*�2��U�^S���;���Q!T?�	�H���J}��Ƴ&<4Wc��8��L!Q���鈨ږ�'�����) 8T�a�����{ۅ���2B��P7��a��,8ˁ?F��d��S֦�V�X��G+V �9D�M���a��U�w��4�?�������,垙n|,�E1`� jm'����2Rd nM
��=#�j�3=WP!L�\��Ss���`�5�G|Zkv���Ğ$�&��oK��y+�܆AH*c7q��(����*S�)���F�3���\tb��D�򯻶�<�*��e�oh�v��F���LoG}��cR�ǎ�M["��j�6��C���c�8L�A�E��
�`��9\�]��_ ���t$����� �(),\�W��K�|p�7,�ɗ�y0:l�n'ʙ��*��r\t{f^49�F�T�����A��j�na�0��m���+��~	��;:)��w�dT¾�z�Wm�������"u�|P���b��⅊1N�����WsO� ��%> ��^����^Y�z��s��+��08)u ^K���z�V/|I���1�����w]��dރ �ԗ��n�=��(�I@d����tfYe2:�#�l���(8{h�R�S�$[@��Ph�y�0�7�e�S驙��c*co{������i���ng�'��>,�L�9
z$�Ͼ]1n��e�,	h�iA���h�7��Ny3���cc׸�t���������u����-0���m���TO�YQ�;�ȆU����倬����u�'�F��PG�L�M(�]�l�|P{�[/�b3N26I]LN'5���G�� ��
ZP+�mދF@m���U< �ǮT;�L 
�pб'!a���,�#P�<��&�J�R�o�Ym��0����������?߲z�M?!Q��N�Q�H��)��vܥ��ڐ\,��p3Y����AU�w�r�珪}��m�w'6��e��}ח�2����d �9rPI���.Rc+䢴�b3}Mɕj�T{�`��f�Y��\]�T�Wh�@e�UN? $���W��u���tw��:ew�?�k�G�ԦH�(��^�[�˖0�B�M�o�6z�F��E��q���:�1y�ҏ����r2~�,=]�[י��Nː�0d�0����г@+B1���)[��RZb��piI�؎䝎���0~VGy���׉k ��&rz�ta��B�谺RG�s���a����P�^��I��5 +��u��N�sJ K�>.*+�VL���w!���9�,jI�#F��F.z��bi��Xx�V�c��*�b��sY.uV �Bxݨ>�*���:�uP�M���`����p�>�H�T����:��\����7k6K�6��4=�f��ͯ�{�r�����������1f��>�w#$��}��l�݅<v ��]tc���PM�l��=X�yP�υDʹ1� y�3x�	p5,+��͑\�l�n\*��C�K��,���HoUV=���:�-�ڴ&����36���-�Þ���	k=�Ɛo�(%%>!c�k�^�)�i����8�-���٘�ho"���Q��E������mFFm���q�z�5��GlNV�mvb����� <5�򴒡;Y&'��/�z���D�*�1,��*oVn��B��#�jaz�.V�A%
%?�ɦ+c.��R*񩻚� Y|e�r����5p��+d�Vu=la!�W���?>��=�щ���[�3ۓ�[7��x��I��-���Ů��%�aՓU7ב�(�</!����=I���J�}��v�-�Q]���G��E���� f��O�-�3i����5�Y��H��5��|��'j[����D>��kt�w,k�G��p|�
ߡ%�]7�����VԶȼ��Z��R�{����r��ߑ2�*
,�W_5_k�J�=�ډ�4\���g|�q
�o��H$��/q�6�qY�N'�Y���׺����w������1a\VúhFQ���1bE��Q � ������sBz���G�"6�RE��Bw��v8�����|T̄���s�[�^2�U�t����) Kb�{�L�d��Ȟ׹ۯ��-�n�8�@�q,��!����0i����7q;��upt�aĀ21���Y����?�h�9q�g��,vk �"�3���v;l`�w�I��Q�=N.�fj�ő�<����&��4�������R�c<:1����e
?�~��s��/&��ц�HO�!t���C/�TE� F}f��H��Ћ�L
�t�T�ힸe�:�U4�miy&+��4k~���!X��jd����x̑�Y�'��e��4�E��kX�н-��s�'�b�%"%�`��` �dYF),ZQ�(@L���GϗR�eUx�CD���RV��T���1���>,�N�� 5����d,�� )~�M��B�8���}h���6ֿ;�Yo���I�T3��#J(�z�7UQ���[��7���P�? -�8�}�����j�@����ad%��[�%vt�n9i\mo�(���'�HR�E*\�m��E͒��M�\%��ǻ?�D+̭zC\f&���۶6�m:�#�`z�pJ�d6͵����tR��"�r��;1��G#�x�=_���^k���Ցm���w���k��ŀ��]+xڄ�'٠d��<ĳ���W-t��IW�a��(�֪���� �kW��/�m�žX�V[N�z&�튾p�&̿j���6G�~U����/�X܃H�`[�Ys��`���O�ƺ�Z=FO3��3�Ufl�?ȹ5�_rF���sN)= ߑZ\P�ъrZ��Om���vE�,�(Х!�;w��X���n��SsL����{=[s8�m,�ź���V[��SV�];�佄3�l�mf�qbt�f�-f����cb�����@��|]��YMj��ڥi��kQ�ؒ;��R��%���������ʭZ��ת�vH�1]�V�h���2�d�^�^��C4m��U��	�j�!�;�g7T������"�b�o�i5ֹ�/ܳ^�� �%�'�8�5�A7\��j�q�\�X�����;�� �D��5X>r[����Z�E�9A���Ȍ���j?��V�|]�k�k�7q{�>�4�N]iަ�y����NS+ �r�#�5@�EJՁ�������F��e%,�J�������@����PQ���'E�zU&����w,�S-��5�c��;�AxP!�a�ӋL���0��k��Z}�J}�����n��+�
�e�=DN�,>e[a�F�/i�7�G�������ݨ�Ap	��c�ߎ�rc���`��?Ѡ�:�ݥ�^2���<�8Q��كmӣ�S���<��W���4 U�~���й�ӧ-� c��y�Z�\��a�Zk�7��qǆ�pG�
(�6��JB����̍��Ȇ,���x�̱$;A��ނ�U�R�wp�2�G��b�\�y�����ӁT��<c-���
�H��]�yPة$���$j�k8�x&C�����aE�&CD��s�a�5"A��wHz������tӁ��DH����K��ڇ��a�h�{���TC���Ѭ4���)�#M��+�&?X+Đ�-sH	Ep"�L<V)���:8�K�q�W$�(<3��ՠs�������6��F��e�qJm��9�	
I!��
�[WF���f�I�QQ/�hF��6�,kg	�Q�$�o�>x�z~,�O�p���W3���(FEӓY0Q��CP�ϧ���p,E���Ó�|������
ZI��2;��G�B$�T=U�]D{�N=�5����ƫ�{O��r�Ԙf�KK<����f_�QQxb)r�)6i���i�k��%+I|��N���M�?���y��eZ��`<M$A��H����5�<���F�v&t�� �-��AO���������Y��kP9w�8���m܁�Rμyz�Բ,-]�K�;���g�6Y�a�Ipy�$ث;��m4��VdK�/��Lr�}ň^SUN��l
J-店H9|j�k�&����h�'͈p(������������`6��ɦ2�C|��3�;��'������F�X� ��)伱��v����n��ۮd�$�s�z�A��2�(�b���x��3���P�tzԙ��ٛG�\ОmI��D���nWf�=0L̬�%�^Y��|9�>Q�VW>�[��#>2��w� �����>�Ɨ���,����1&�����zΧ_�k}i�
9${7���#����쥒�O��Tʜ,>
��,�����`�yz� ����G��Q|N<j�?�V�>��������������Α����fb��Aؓ�aN��Z���������+��I��v��x�qS�P82"{��^,��߾5_J]2K8]fQ���)��`~������F7��F�G��s�k>B�j3V��J��hH��s_��G�|���@�VC��̘���}ϸ����pQ��|�=�Q��ړ��+
��`L��΋�+�e��v/�d��L��l j�.	#0�Du�|�F��-Őe\Z�J���k(�����k�F�K����4\��)�L��E�����+gh��ބ��WUӲXB9�z���տb���4��=a�<��e��p �ը�	�,��h �_]�qc���[6@%(�B�Ar�%��|���n=ޯ�(�m�W@H�P�FLa�E��a�o�N6pJf��k�E�� ��	��ܞ�`� �a����1�ڐ�Z1
�	q!��_���L:�ť��/� j�M��9#$x���3Mi��}�u�R�A�����=�b���f���8���iE�v*��Ȅ1Nk�%'��W��Nڋ񎻳6��bp�k߄x����{�R'�z�]��ā�m���8��.�����y'���dH�}�/�c�%m�J9���-U�t1��Kw�z67	�Hc[���Q���R�Eu&�r��N�PU�g0����s�6������쌼���j���іTi�׹����E�r������qu�8�_� 7�|��;��]����w��а���-�@|9�4=�a�ۙ�)��r�=uP{XT��@z8�6z	PEY
M�-:�R�Bo���i��������Ƒ4R�	�
�2$�mя칫Tz8;�����q>m5AΛ�$\�;"۸�_��L�,�7
�T���1�|v�����r��w�vϣ'*ڷ��|�gQQaF9O��-����0[��\�l߰��R*�JP�4^=�l��7@�5�3�>��I�ww�c�z�k�F;7��Ǩ)��Z�a˪�]S�� �7ǁ8�E�˴�:�oㅫ���5������ ���H�hS��| ��J*E���~���
���S�Rj�8R��򣃪!�!�PG�:?�WF9u4v �4.r�[�;��N����8ق��4p&
!�.o�^�&۴2�Xt'RU!{�a�Sj���9���lc�t�����?f��`%Ͽf�&�x,	ԛ�P�I�竭ֈPTJ[c�J�<���,�7����6�&y�V!��h/ �P����>�7闸_�E,�7c�$������ �8�$�"���cܙ!��~���!j'�2�4�(��s_�asTJd��%չ_�	��Rs�q��/yZY���k�?�M���d�v4*�?� J��k+�����Ӑ�jjlBN^�� �݀�]�&��ׇx��կ�k���G{ʜ�=b�r���G`���\�;��ߔ��2�<[w����SM�:,�ޔ�i?:���G�5�k�1;��ܣ\%�b��naW���������`��`�)O7��}�L?d9�s���m�� O���r�:Ρ�x�4��])v,x���]i��$�5ۅ���a����Cy(k�6V'�iTl�b�f,��;�goY�~"�볎?;��i�eeD��J�^j���r�����$�X�C]�a)�,��,�&�SS���1'�q^�O` mկ���*��v��84�=��Y~I��Y�����.��l������L�I/4�66+��ܷ��(K�yߛ3�O�����vZ�.7�O�\Q4�����Z\�q�+�C&��W��=��I7�A���'*����h�(��#�O�Y��T��o~����� Nժܔ6��B �^�q^�n��F�>z
��U�rlmF1e*��g�&�� �����J�v�=��*Y��$XA�0,�a��q�Y=3�Hs�ُw�_�V�)Ew�bg ��.	^����i,�/�7*׸jJ���@;j���_�j4:�h��\ޛ����qB��i�9��֞�=ԓ�xB���6b'����eNt]Z-j�0j���d���4�E;�V�o�B2']��	J���.���w�F�M��'u�C�'���z��k7#|�&�1V�w����})M�@����f�ER���/M�-�x��e���A^;|��-o?����N�/��!@��:a���y#���t�����w��s~�Z��/V�2�����}�GD�t�^�e͐�>��_�Y�λ���Ǒ����ʼ&�ǆ����%�[2�����X�����^{N�F�����k"W�P����.�&�\.�C��(Է��+���uԬEi�1����]�����~Q���/O<�%8���G�����xN�X8��Yv�?�3��P{���-�!���r�Ľ�=�|8��?��N�^+��05H���[{���	�U����aR����������m|��fF=ނ�x�'�Ռ���\�X�"xr�#x�Xh�2C����:�A�q�<�gK7�6�0�����oD������3��Y��j
��|p.%h!�~����v/b�<9q��q0�c�g �l7���y������q���J��EB�=б��A��E�?	�"A�ѕ�cn����d^�����.�*���3�T�'�ܺB�q�"���CD[`�)��u��=}��/UE|R���G�G-�ྥP&�h/��\G�)l���X����X�57�<~+������|R��Pe�p�M~#��fYr�o1L�>
m�j	��F��������<�U��O1D�>�I������g�[Aǈ��36�L�y�P�#��9j?H՗���G��i��[��o��x�gË ����Dq0�@� t��/)p�x,)|j?}IYa�7���&
SrksB�'�s�w�s��t�
�%�� q�hr<_;�q6�pN7Č�"�w#Y5�!Y�8幝�k�b]�>S��A��,D�m��=�_i�p��1ǣ� ��������$�c�^���D.S�ڇ=e�z?��8L1	�F����O�h'�9�@�4��(�Ó�d�T ��ه}�ٺoWt��&�|��;
+�%�F}�+�D����eaX�Qr7�޵rY����P$��U���T�OƲH �<�ԡ+A]�!����ւ1�ب՗0���{Z �s%�H�R
�-�����,��$��|��Wr���/���	o�S$�+��rW�~��_ ��O�]�oؤj١�g������a�)���*�)���u�BTK�3�>>~�6�t��D'JR�oŲ�dan�f��祧��'�r(�C��.�
\u$Oi����v�O��.բ�Y�:���\��s�]��������Ec�g.�v'ծ�Q�-6�\(BB'v�A������e-?D��L��A��M��L��#(�Iz᥆@���dY���w�\΂oǈ>���\��(Qp�0�2�����Z�5��j� {�AvF���3K ekh<7$��X��b̝���:3�3�U#W�r���η��D�\��fX��*�gX��Uf�0���)��TV�M�^�4r{ϼ��WJs_r��4���$�Y�,���&;���t��1Z�����iK�i6�4����IW5���D�|^���р8�[��k����X��0Pxw$U�Dh ������D��cH��<�u�	R���fϸ;�@��9�h�����5i	/��~��%���g�75qǽ�j���UL�'5Ry����5���B�A�År���M�K�n��j�{=
��"�C�^�����"G����vt��9��8ol���`A�-�C�F I|�L�]��/�ϩ�����\�%�������*A-_��+���i<�߂�EB���[�w���^ۡ�dI�?M0E�"����m/�PY�8-�B:���c����l=�>e2��^��W;�E�4we^��|�f�[��\��Ρ������c�s�G���a����(%��n1B!y�8�!��#(nE��Z���m�6�Z��w�8~
������QCN�\�Bf]����	2��Nl8�*�Z�	s���{7G�Z��!S5������4�u�
�>o}�K�>�8��Nu~�?cT���y���0e����3� �5ڪ���2�A��ϐ���p��]�Ij�B �օ�<�BI���FO��p$�v1��Z��m��o3��0)���bw�V�$�*�^�-�����q�S�v����Y�{�/yw+�d��]ن�!��^G ��i��D�Z��B����7�-i�ٯ���Kӟ�6�'|?���T�.g,
��jR&'+��w�_�g��̚K����Z���ZaW.������6| �^m�+.���mC���vu{�[b�pa��o��v��U�G�T��H��w�[�"G��"���z- �Ҍ�i��wS2�$#ҵ���������;Q[Y8X�R���y��S?�L�t�n���x����N�#(zw�T+�"T`����8I����%tY+������м+���`���ٴ�����:)&�Oa$ڂ�8��s����U'a�y�{U��ė�vJ�<J��ɟk���N.�' Ib�����W�p}L> �
�j�?�);*�2O8���{#�k?G]j/��	z��u_�*�],�#�Qm_J�D���TI}�l��V/��(qjI��
S�R�٘[�� �ʀ�_��C��M���+n2z_FV8B�zX��V���� _R~z�w<>^R��G�u�b~zٓL�
���}�h͋A������U�tb���ϣK��G�Ԥ�nSrW�Q��	8�!7'�n+��Dr��`��7����#��n�]����:����@�LC�%
wT���K#�L&N�w��fI.�;���#�|�z�Z����͏�L-��ܓ�z����RH]$�݀��/;a��O�ګ�d��e
� ����S=Ax,<-�e�{��>c&�o� �� �·���\b�E�*�p������y�H(D#�v�9���A�e�f�� oA�����p \���]�#z,�������x�Jx�j��J~n�DX��N�@%؍C�@��1s��i��+V�1J�X� �-})�P�+��x��]�i�iL2Q�3���ٳ�9��[G�ri��w06>>��0 �b�3�!
/0��A�a�x��֓��9qf��A�|����	��+c�	�<�l<]yri��M�?� ��ܘ+�!"-	�ps�oV2�Z�bP�7C�f�"j�;�>=��0��9���6�c����y��
oJ��.o�Uߋ$�V��\���栖3R�TY�#%1�b
�S��,v������2+GSX�=���g2n�E9>�.��טp��׿�Dᝉ��Z���kqߚR�g}��z��P�%Nl���X̳.<�,���;y)Wc�?��N(�gE��������G^i�ixX��<20z��񾙧����H����"�S�!�/���GD�eQ�By;��0��2�t��j�J,_H��D>�*&��e���YFfX\�4Z#�6�4f>!Pb�q�R�%	9���s���%�-*���������5�����6�CP��� ��|��=rD9V�I��C���#�N���I�d��(�8O)o��q)�C��t	&�!�W�ny|�j�I��d�r�D�e������s%Vc�t��!8_ �*��\ІuJ�%�\��^�:��d��^PVu�90,m͖�L�K�\�9�`�2��;Xm�r�6H��ΪD�k�):��%�h㩉��`W�6��僛GM$0�J4�+�#m�JD��">7�ц���؅<��1�ψ�*,�0_��9i�3�("�\��G��9Y��:�ś˞K��q(�Q�5˝�$Y�j���3��#��arzD�'�}W����ʶ�N4��¼ǃ��Kr)A\iQX����c�Hm��ۢz�ΆgnX�@��+q�(��2q�o7�ۤ�L��f��@~C�{{�aY����85��S��M	�%����\�*Ir�J��}����.��5��@�*�'��(�W�*�be1����k�����|!"�L�dh��q�a3��(>�-���D;�L�n ���^���ٍ��)���Gp��c`���o���'8L�w�{Q�h�$����X�E���d�o�����B!��,6���_��#u�D�BNR�m'�ssLōiU�Y�������+�_���p[	��-	͠4�^	=P��31�K<-���o��0�lBe?�R�˸Y fm��Q�jIi&-�A'F	�Z�$=u|ρLT�Ɔ5���%YΦ<�Lp(�/�"P�qS�J���ށR��U��j���y��(�]vڻ6�ܶ�A�f�����JRb�\��K���P�P1�G���� ��F���C�K��ݹg��ĬnÍcX��]�H����f\~��X3_��ۜ[�W�n�Ώ�l~T#����+�ƣ$�g
��Nd�H#Q�E�;�|���r��u
{9�^�"!٦۵bh��z�Z�W���!Z�[
���́�m#�����G)\��l�B��O1i��6B�V��IG���~���g#Jb�0��vˋAq)0j����;�0�O�+]i��.j'�R3�5~��T���$��s�����v\<�c~	[0v�������Qj���=�w��ɵ�0w���Iܻ V#��RH�;�Ѷ�� �c��������MK���F=����ƆťR���ry�lQ@n�Ɏy<{��)�Z� ?��	��jz�ީ���S���HV6�LȦƆ<���>����gm��y>��d��:�;{��U����qF42�'��1�`�[�.�I�����l&�U�u2%�呴Z\K�8�-2���T�X�l�����[�M�d~foOcG����]%0H{��o ��m��ǖ���}�S��M`��1�t�E;V�K8"f�&n��v-�xY���ٜ��mn�,2l���~��z�S�<��^y�FmO_n��C��=4��`J�/��P�<q	���W]�;�r��9��9���y�g�'z��A�y��X�ʗ�N�����WY����@1��v?,;p�.�FN��xB�VX���&�b�c�pc���ge3 '�'����$�Bs3���A1����q��	�}%��t�[������!P���^mk ܓyf�9�?�F��)s��_Bt�.��6Z��!)�t��|��V������W�������EB��N=3m��_ ��{4Ҋ��G(�@~�ȑ�����)��~��ѫ5��R�87T�k16�������f��Io%�g��z��3��*��J�5X�{�Ξń#�0�C̯G/��$���]������<��MOf�܌;'�Ó		�龨�}�j�|�mi*uC�������#<A���:#+s�3Q�?x�;Pg�ǩ���e�L�ρjbv���A�8��3�H�������Y�-��>�4[��w~y:DX���4�`Ŧ��~���SC%���1?��w�\�#�%��#���ʠ����U��P��Q��PSюק�����i����FY�|��du�6w
u�_W�����76��HD��E�}��F�Z4V.O�|�Y������u�ZcX�N
��������Ԫ6�_���}�ǳ�SG�Z�`��n�6���O�Y��9T!��
K�/Â��-����W^q��|k7ؕ8b��Un�t�צwH�Qq�JA�,9�?����"h��d�x)j�l�xR�.�yo.��7�R�	���3E��Q.8�edu7-��*����ED.��Naԣ�>�T��Kq�Gia3�v����OXQ�[9��=�ҧ)����x�RF'ߕ��t0MZҙՋ����� ݁s<���},W��M�_�a:(����)W�K�������A��5�kz�T6�)����>��[�_)�����nAfd��U)&L-0����]\$���ˌyO<�sAL�k3܇o�a��}^�{ ~v��oCF���,9O�H�6�d �/�f�B!�R�1hw���#�)r���Sf����P�P��9T�IZ4_H�?IH��Ҩ;��m&�ߎ��/߼�&�k�jYk�qH@6�5Z
V���'b�qH����M?pc�@��Uܿ�J�:���F̺�l���L��:m�6�G��>��Hgr��~TǷ��
6��4�/��[m$OrKm�?iwO{�5-(�<^N��HQx��]��%~ݤ��*u�tY�|#,Z��ؐ��}���o_Ψ�R'1���B��� {'�P��-,���O��U���q#�k�}d,%�-�ѹ��G�0h҇��EL\;��L P��r�ō^�p.^������f�tO�Y�
�L��,�I|���8��b:�w�w,"��ڟKE�d�J�9�m�g��ާ����t�"�XurE�
B\[���JY��eӏǠ���BQ[��*�l0��BɶY�Z��p����mYw��]����[�z>���6rXnJS����0���kCߊ룾uQ���Wz����W�s3M�;�lK%0�`_���%n�)��� ,��ǪD�ж����v�H����V�_��d�A=��7�9���Ō-o��U�_<��G�P�i�bp�0��[�¾���}���C�U�7:]C�'��2ᄖy;S��(�B
O��=C���d����g���hu���X���:<I��&��?݋��L��9�^ԅ��4���E� @�+��7��	'��A�kK�1Zjm�t���L��;uR�zq&�z@��7�("p�c�ê_�xk������(�^�	j�����������8G������Z���+Ҭ��.�y����Vi64�5�ST&<�� �YVQ^!é���LKh~MO��l�x}�	mvA%3�V�:c=dC�*�*����Nl����{��x �F��Q0������ߚ0�O"�J*K00��A�� �H1��Ѫ1{���I��9V�O Ƴ�Li��t�L�(�|$��NF�N�Ҡo�7�0a}Si�s6Ԩ���o����TU���x��Gx$�B|��#���.,��V"��;$�tUȌth��4�=XjY͠A��tJ��aO��:�#B����Gv�s�T;`@�@-��h��΄撛�`F@@�B���^�>������K����O�1����Ma=8�����T-\Ә3����,�,
 �oJ��s�I4�8�a:9U�K���o��b�o��v���2�~�p�~���eT�se(J���؇�����@����k��!sT�cb�[�3��.M�@�\zj�O_�H�>�������@��|1z���pq"���:�g|c���g���FZ7*�7�����:��e��c����U]�ʴ�L�<�D�J�@����ީ��,CT�娃�JYW\�ݠ#�K�[AU�aa���4��j��ڤAjN.��ݶ`����m�{�Z�`���@a>[�Ѭ,�s��thm��vDb���u<�i������K����.�p��}� K!�J��B��`�qp�Z5��0���Q�"��<�&�ፏ�;�o ��x�m]E~ԍ�j��N�n�˝��B�+V�e���Dl+�A&S�����*�7̱����,�������Y�<�zV����&Bٖ�n���T���2��
J1Xk7�c��2�����A���.[��XOZƴ	�I��!����0\��I��� RH'A��);��G��&XW��l�,[o�c�Z�5s����mSOm��,aݼ&��)j2m
jnRR��r29��;�t��%D���KQS�[y��302e�_��*�r+6�� Z�e��|�p�\%D���`,vcЏ>�pE<T��=2�X�T��?K��7�9Ԙ�sb��D��d������	��w�����=cv؞���Ũ��h��.�~�丶�=�QZ*Ʀ���7W�� �5�^B��Pȷu��W��i'*���Ѻ��W�f4��㉶�����ڧ��"V<I#Ii��ߨ�ƍ�8��Fz w���3w�9�����ɩ�7Q��B4-R"���V��H���+}����Z�ĩ[�#׻�6d���ο&��q���N)��]���QWa��<;����o��&l����9���g %��[EE���(�L��+!�����A��� ;��Ō�c��O��yʷa}��	�\3"�����O��Ũ�hG("#H�{���3{I?��p��&��������ʠP8��	bN1Fvt0��Z1ʷ鳮��u7��(�x�l?Eed5�$>�)���*Q�3��Yu+�ɒ����qj��[ͼ����ݦU�˞/��a21$�%/_� �����2T3�O���M� ?W�~�/�����_�N��i�[�(���^ܛqT��N�^S=�u{��.X�e*���.�b��S,a��"�Vk)�P�4��ɴ�]1A� C�j���X��#6Q}(���ˏg"���eU�</f�̒;����r���_�="+�v�{�lV���p-}}{�a���yς�K��P���]d�j~���w���R�Q��o�QĖ3�`.���P�^�T�O�t��j��\Q�R����'���dZ���),1��^(H����̭��+�Β�S�Kx��6������U�c���_Op;�:B
�&�Qf`&��:$��F��J�Z4�*j/=NC"ge����I>�P��a�Oy�>�����NJ���^����z��|��!Z"][�'�Ѿ��g��H(���O�(���E������/�
��͞f~ǲ�4c���/%�-FҶ�\p��R?��@�x�zU�����&����Y߂}A�`�)UHځY,=�>�^7ris8�Ci������&�0� ��*�)������XN�h��lPt�s?� �&rgD����꒝��Hl]]���,��Z_5b�*�f�����q�ø�s�����^��Te%��s�sl{V��E^���I�b��{k��e��M+����Q\U*ˇ+ۛ*�j|"Y��r��5�i.��9�2OV���y�\�b�n�8�@�+O#JSS�ϋ�{�$�J���j��9\�*�� -Jm�2t7@�K�9�T�wZ)ٻ�P�+�mL���)�a<�2ώ�P�\T��\��zM�P��{8��	G���ٺ/p6��?(�h!�#	�J�ң��tM�{��=GY?�!L���?��wȧ���A���۔���J�6�@G��r��fda=};.����@����������d��Ƥ  5���'~�z67~&J�u���QJ"�.?����0����p2�j���#�xQ|W��}�e+H�X	�U�z��Є0�V��$�@V�=��!`�R*(�m��~����s�;��t�6I��j�Sn��R��1����Zl��N��]�!v�����||�A�&�A|s_����b���	��������`��ՋF�`�#��z�h�5'�0JA=����L���bz��q��	�z,˄�Q�l$'/�j�w����J�Q��>(��P���z�d�F/H��HOp��.E� <��q,oی���ET�u�Sb��*/6�C�W�)w�� �v�Q5�&�z7A
V���u�B�����yo4�;�u�� ��bӝ�˯�vhg�p\ul��)��<Ni#

Q@�-QC5���(b�F��b*,�j�� >�����A1uNyt.x٧�A(+��Oa /�����B2���@��'	'��De�-��&����j�<~Yoc��R��o�s"q��W'���!��l�>��j�N��8?靍����T�Fͤ�w�G�r�T|^�D��{ȷ��Z~!08&��R�]��� �P� ғ(����\{���*O��P�g4v5!�q�T�s�d<ܼ�]��N~�o>��<f2�6!E騡WQ	ħ��z,Ĵ�����Ո�[�m�P�"�G���G]AxY&��h��?I�au*SB���S�u�v��43 a|��{u�M��ݺ ٤Mؙ������Y����ѱ�n�nQ��*a�ҦmL�5tU&�H�ӥ&��.��G��톮{	�g�6����u��ۈ��6���}�y�W~_�+@ǽ@)��rW큋ݷ��&l�
n&�4>���4._j�u�ݼ�ѫ�$�x��e������|���$Nٳ�Z�Vˏ>Cm��T6�V�f=w�鋗��[�y@P�&A��8�O���,���u6 ��?�v�	@jˊ���5	�I�/� ��$N67����8�V3 �)=��d�aܨ���kȰcN~
?b�މ'���ϔ)I���K��_�Mk�d{c�(9�-+����m�<ʊ��g��k�H��U�MИM�]]^!�XZ�ڞl[����{��Ǡ;��1ga�	���;�O�ڸp��v�:"p1���L5s�U��2S����!�*}���D��Z���B��� ���9ׂ�vάq�1O�o]DMm0$���)ű��1��}�#����Y|������]�LYi�M�Nk��ҽ������	bddςs���H*��K��r�۩"��
�m��5(-1��jw^G����b��IJ��[����X� 	&3��y)#��5x�u��6����f�^aaW��L����~	7�il�H0j�;ȱ"�K����(���W�,�fm�R�V���q��Η�uW�_]����@5kJ�0j4���҂LF�FD�;L��[9ɭ^'HZv�o�y���:0%�*�o�\�2k�g�SJ��	CJou����
,��R��@ z�q0y�a�¬�b7Xȕ��z���S���C�UuR�G;��ӀEVq��Ssw�,�T9j9~�s9�֎EO*����mP#`��:�˛����\�9U�|i�� dck�`n_���!G���i�Tg*ij[��A���{&�]��#�u.�[�Wcl1/S�E	�(�s�G�?8a 7N��0K���BQH�c.�a�w�;�����D��U=�E%'O����2���I�D4�#������W_q9c�X�yr���4�z�Ŝ{�5VZ�	�̲	WL�8{g��� ����X
pvPn�%X�d�z�B3Z�ZN�%Y���c�)��j�U�-�p9/���t�G�!|Œy�/��R�|���\���ScAԶgH�X��d�%�p��7���p����B��\૔����������d��$f>�+z�f�Q]<k�2�Jfd�&R<��7M#OpϘ7D�T��aR�Vܼ�ZJz�_���d�e�!K`�	j ���3�i��i��&@��My)�,�ۑZqy�k����g�����X�H��Č�)"B�_�}�_����F8ϊ����g�F3?F�4F6�_��_`���vEJ�k���
��b�L{+�²����E��Bh���mBc�m�[O�+2�Ϥ��=��h�������cع��G�:%y`UP��K�5w��(����{��@C����l$v�O�X����j-}ߙ	�|�-�~?�LP@VT�.d������{#�G��t��xР���P�_�PP�e��Z²�p%I3�^���M���
؊�K<�
u��U�B5���"�>�K��/o��f�l&*��(<2���4C+��롛�~pV�%��1sY@}U��^��I��cg-�>�/�YdP�uqD�@����jB���G��E�C)V��	�_^W�z������xq�"��Y輺?�N��U����U|m��p������4��r%lz�;�[Ӝ�
s�"}��`�g�;U�nE9�ˎ�Yu����1�EI�����0�>aq��ן�
���<�6�� 0/*O#�Ib�!��E�ßh��ؚ2M�	L�OG�vg࿤CXU�p8��T>��;��L�&�������8�}C��3zR�b� 펳���)��B��9�q5\�P�`�rR�g�º��7�=��D�X�5�Q8[E�B6l+���Q��Y��F�v�� ���,���4��z#��2���P�êӔ�vV����Ӟ��w�J����'��뫣ι�G�Z�� �C+���-�dS���?`�l}:TY�ټ]������,���Z����Qp0�kX�ٱ�ک�}�U� A���n�p���1Ϻ�lm��p|+��1��N#ɰEr�+F��Rbv���X����c��h
��h��@#3�9�; ;�5apr�]�2�X'уY4���-�$b�uJ�Ū�L���B�����Fj:[a���S�F���A�KD������䩠8��Fu����X{��ǀ�V��^8{D_�tݛ�th*���&�6X�3Ѩ�^Y�u;b�*��lk�ߗ�̜���>1�b�2\�cK�6��=4H��9�����c���S���|8�U��J�z����� W�S�ɿ�!�L��ye�&�_ R�2�	:`-��0�^P؃/��h�:G���Ke�M-+�E�]�H{c|VrB&�.��_Q��x����P�cl�8��R�'f�ߥ��eеO�M�]H�%�Ms�w�U�FW��pl�r�-�ҥTD]�}�> ��Dߗ;�m}�_�(����!�k@�Zn=���3=�s9w#����/�=���h�3h_R9A����'J������1v�}�*�����kH	�9�>2���9�y��G ����IĪ�jMs>�b�0m.+hѺ]#��Ķ4��BX����H&Ki3�.��P9f��'W%	�\��$���t�N�6�|�s6�����*e@�h�Y"ӥ�� �ۯ؛���S��l��L��SI���o*"z�
N/�����W��������5���"S�X�J�	(<'v*l����ߖ:p��S���3�!��N�o���8���ɪ�`#ǏT=
��S;q��,ݓ���oxn=�Q=U9��DnK���MtRo<��)(�~&(K�5�-Z-��QV]/���d��W�(ߧ����2�G��FS�[�e�z�9y%%����G�k���&xN.���W⤛�?����TG�Aޔ�f�|^ͣ-��F6s��~����7�}(��1��|C��GC\���<��s�Am���܏u��3eVl��zx�{�Ru�D	w�G��?�A���:(�9c��2� �P�{�߆�jt��%��A�q��5�T(��ݭ�Y)����Ƒ�u���*ԑ.z{���n���MAG���=� �b8f�u;�R�$D
��w5�n����`�7Tf�T��m:�H��up�N�Pʓ�[�d�w�n��Րڅބon����Ml
xs�ЀF���~v���ǯ,q.F��P�@3b?�X#�(;=�zY	R�׈��͙]Q3:��户��	,�|(#)��1��f=p���|Y-�I��\�p!�B#A�����Lqߡ�*� �[�a��ۙ�y��c����m$3j�n��;f�C������@��Yg���$'
�Fh���W���h��/~F|@ѕ*a��$km�d����i/���rj�`%�gn�F@�����n1|���	_%��-��7:�T�#���8�[͐��O��/�V����DMa�47,oJ�"`ƁE	�qԛj���L�*1N��� ����n�"��R&�)��um0�aAyj���	p��f���x���u��a��']� ��lI6.wlFS��G�mdi��O�n����-07N%}�\��hz\�ޑn�`T����?S)�ؙ T�Z�.`��As��.V[\� �����1p)�g�SYc�R�x0N�3I���z |� 2�7���mpM1)��A�Y.c���A��v���#��"���fH �[�����]�����n	a�ā�J#���lWi~�Aw��	�C���m�F���èK��s}}�{�2w�����f�,ꕤ&�X�{��k�W����b�W���V��V��BMdG�{ �v3��б��х[����"���PKճP� ݜA��6���Ղ@�����l�8����|?�|�@����Mq��D7	��ۛ�"�B-�=�G��:�"o��
����`��G�Q�B����y8)H]AB��ú�e��&'�r�.��w�b��ͤ�G���Մ����G9R�(�9�g�X���5�Wb�#�BG���B@ɞk��ص�т�Ht��W����L �:QQ��9!	�_qcr���aC���+?sk�z��DPJ����S3y��(�S��+ ?����;���OfGȢ�#�Ys}td����TÎkL�2��EN�Y������A�9Y��\[���$a߁�����N�YB��,aLk#���KFA>$}{R][�4��H�L�K�����f�^X�T����ߵGV������O���hx�M�E��c��)aX�4.6A�*��1����|T5ō���""�r���9
=���)��tG��MwmX8Q0��;C�{|�C�!8��t#��3Sτ��	}� 6��*�2���ǭϛ��!%�� �
�!:V7�V�Wvx�B�����E��}�1��riگ5i�����	a.�&�ɣc�t��P����*_���-���	����$�z��ۆ �rFb�;��w)��M�e]����D��բ���O�8��Q
{��1ӱ�E3��`2R�<L�;�Tٍ[h;���;�_����^3����o��W.1��S)�P��ӗ4'��W?훱�A/�2������c]�r_Jd�y�L����j�{Q'>=(Ɇ�\�/0���Y��p���$���ŉ����n�1�g�݇�lT��9|�4�rY�4q��}���U�ć�i3�m"p�'רM��q�q��Ƀ��	��f�MúE�=��c�e���S# rYy!�U�����-�Fy�8{�O����w9-�n�K����)c�ɱ��(�8��%�mHhZs�1�l��ġtz�ew��W���0��p����.-��Ƈ��֌��v��\���{�E�T�$��}[����O�h���ΩԄ}����!d����N`���G�-�������Ƃ�9�?�b��ʄg�)�1�9T���O�%��Se���v�H?�>�vW����֜�ܩcm�����&W٭�iE���k�d&��i���Y�I��KT��w�+R}�.�T
��
��ł�8�So�Ǚ����̂��!�c8v��p��jV�I.e8��Q�f!\�%����cl��sM��o�����v ��}=��bp{�ˣQ�Z�s?D���(닜7<t�b�	�̈_�J&�T�p� �mv0u0r	V�B)e=:�d��&�������M"k�*'��
a�%�O2�A4���K�7���@qd����r;a6ȝ����"M=�ԁ�E<"�3�.'����L|�w2�W;���gN��$�5�?��\-���*̝�F=�5#ߧ��㪽N��!�d�g;L5��q'�ﮖ��4�pB�'�5�p"UZ:�&M/���[.�j-���­����c�%���pQ�]r�g.��������%Vс�����K�C����	�+��&?:��N]�&���>rXK��$<�!�&*������+^[p�7�=�0�L�uQ���Wy��<� bj�Er�L�=IX �L���ؼ��,\��<!N�?��Ɠ���}&�U$6��G�N��^�m��o� �y�ɰjֿ�rEA���Y��p��]gC���fQ�,�:7�r�����y=�X1�o ht�+�SI�v���#�5ɴ&Ƴ'���eT]n"S�70x[ֽ	��Z	�	!ef���'�[��f���T��%���w�`��H�~���-_�D��+�*:&g�ls�\�]�N�ɑ�M����kN0ѓ�_L
SB��`P��X�G���O�8ҝ��^��ߏ�AE��v�vΏ)��r��h�"����
S�ى����ylowY�<��ˋN�����MX�<r�Jg�B�x*��A���^#���d��불�{�I��sz��sd��J�?�0#���M��e�'�����b�Q�ʪ5�w��T^�x7����(l.س���e�V��3�L|Ŗ8�t�p4���E����ᛤuST`�uL�;Ⱥ^A��*[6�}y\�P�ʔd��Qѧb&�q�*���2B�ԁ�ֻ�0U2SWq�-�����7Z�s8��c�1���1I�VG���pF��4p�WWʙ��.H����Q��l<��Ԡt���՚�6k^�MAwYt ���&�p'���?=K�my+V��r���l�)��׍�G03�9��9lɘ��-=�jf��L�yg 9���0����I�Z��ru���WR�M8%��M�7�L���k��}�[��N�=5��F�z�I��~�[�+��׀ !:#�S���C��Ac�⃭��;�a�^�_����ˎz�U���e74���N�)�xjDU;۸�f�y��Rk������#섙�B��#�h���� UJ0V�I��� iUV�iXJ����I���]�ղ���Z0�F��O�`�������pG��6��J?C�rD�����P{����a�(�,B;��y��u��q#4��6V������*��f�vK���<�C�U�bx�I �K�#��|��h4v��-��Ҡ*��G0�*jD
��e�mE��|��up�g8S��F:����sh� ��S|msi�U���J%�:2��Z=	+���Xb���9&�������#E�a4��m�#i�XY��n�[!�틘4>+nфo�Ao>w��x��:�6viG$N�kb2���}���M= A��P���P�neQ�>E[@ty�=��ơ1z����3&k�*�1������F]����6!��z`�Õ���,9N�Ԏ�
@woQs	i��(�)��^�g�]�v�,�F���{���}��6!���ޙ����{5�8���Da)?��&��������}��#u��!4�������E�~���B�
������D�R�G�Dga�d�'{��T�蒚����*=i��18��"���1Y]�g���j�H�7'q�W��Qj�R�$�j0�����(qHڕ��Q^t��嵚������}S�S3�r��|�O�sG=O}}��?[D9�g���l�5����6e��<W�����d'1CO�����!�t����_OFL'*�L����%{��\#�m�0�3�66�����@/J���0o^�1��D����^P0�Q'+ߨ�rD�g�'�sr�B�8�Zݞ��'BK_���#�t4��-6����Am)�sCע5C*��B�8���&,���[G�e}^����K��4{�i}J*�qU�i�a}�����9���Oޖ&m�E/\>�Y
6��&��Az�v��V�c��e�e�G���/b��W��WG�� �������D�{oc�.0"х4��G)�%�-#\]3���[�'W|�D_�(*a��G-�a|���L҉�3���"�s�p+z��l,���Eb����ǧ�c�)�rE�p�<m���.-�g>�u3N�)��B̤C�!�ٌ��3����~��� � �_7�_��M4��2�/
ƛК�@�Y�sd}��}�p��P����(��P�/�4W5��%��O��ad!�z�s�|M�gm$Ã%��D��=<���j�}� �iS�d�H���[�p���$��sV�J�M�00J�6mƾ��\�]'�1{���JZ[��)��O�i����n&&LJ/,��Y���]3r��Uj�)�RKQ��ux��J�x����X��d"� V�e|��3��-\��X��|g	l��4�e^pi�W�UV(K�+A�5-�|a��n�	�Sm=LwL�\)]Q2����	`cl�%��z�&>6��ЬY���f� �Y4�pOu���8@�X,���Z����N�M�}�8෠X�������4:�=�A5��x�G���1��؟u<�xs�B���7QB������V�A.��\._}��0�~��Go�s�(-݃��V4.�{������[��^Y�M^��N�}�xŅ�[{�J����TF�s7��ƁV���1�3�����*�0X�#�R�� ۝�V�۞�}9e3s��6��:����	�2��&Irp����>K��r�k'jE�\��\�)��@�k;^�(Ϡ�a�~�e,�Ѹv�;J� ��X���f߃��L�����w���������F�K^4M�����M�V<�TQAL6\+����� 1ۚ{�=��կ[|��\Ж�"ȸ"1$RS�V��g��Z�`���m���X-_���F۸ue
�ݺ����������lF��Zq�v��j��a����6�N�3�Ȝ��f�������B&�_gDg�zl-�fm�SׇB�b,��:c�n�y�_> �I �pS��hg�W᧗��Vi�k��
��j<hϜ}��q�Nب�����h��V�_Dr�޷̶@��/Qg�B�!}4O�c��`f�����G�D���7W)��aH_6-��+��_c��_~fn�o7��PSBӗ�"ݥcpB"���c���`��.~��i���}9^��'�O�I2��
�O�բG���6����-�-��	�c�`ó�[Ul����n��(i�=� �:q�������S*��d� ؚ�Wx����U6�.�duڟZ�M�.{�͌Ɏ��#�����G%�v�i"Z7o�Y���V(�Fqv�C�9���u�R�7���D�,eׄa&T	^z��*��.�\���HHL��rb<=�ٗ>Q��-*�*~�r�v/��}h�>��Jx;~T�-,���Q�� ���.z�@��e�i8�����������U��ɿ�t(�Ո*�ȯ� �=(��J��l�_��:Ml|�e_o��ZGQ\�C�E*�'��7g�=���x�?�Y,1dL��`���*��Ì+��_hL�H�$�兗ŋf��ɪ���Z�2�2���L �QТ�5���!�?�<1���s��[����s,���M��cĶO���� 4��?�{��]��D*�W�)�:ܹ6-D��I����8�GU����[4�i�t�S��������F�_uˋ}�~���Fm4py���h�6�c\&9�7���){,[?f��M��O���}Z�m���|�=�����#n�����㕉��AO,��h���"�Y��-��^���~o���@���:�`ۛ�����@6���r�~�§/�설So,)	'�b�9Y��mσE�x�Z�����Ϡ�r�*��x��m��Q9ѐ]ƭ��2>��n�|7+ÿ3�Zoa�����rc¸�� vR�b�C�s�����߾�u`�r0N7,��q�kһTƏƙ'�k���Y7�����e���|v#y�������aolK��@K B�47۔w!-�?Ovrm3n��'fH��|3_$71���$^i�]�JYG]����X3@b�+oM�%n�W�����&���w�t�����,��
�����G+�2�@|A:���k����G�(��4�	$�;�-�ϡ��So��h��)����̐K�52x�T�S�'iÖ�e�&���>[ғ��5�����f~��B^*�1��O�z�}�� ��MmQ�{��W�k�:!ǘZ)�9�N h��*\�"$᪊iHpi��X�#y����xf���������ҔDq�+�[�o]����2�q[8.�K��B���l����`�L�;hL^�VD�5g;��Y�r7�o�����!f���� l]��dm�ݪ_���Y^����h VE�G�k�I�r����#�L5�ZA��b�M��u0:�g�	?�+M��t�7׿��u'Gi���|a����g��BxP�:R:sG1)���ZU��b���U�p��x�t�j�#.\�����\l� Nfy��]Ѓ��4'�ƚ�k��N}>$�yQRE_�O��ﭢ�n��� Im�t��LG:�ݺq9 #���J,��=u��b!�Nvw�ﯝ����n�HM�#@�v2�ML���6s��a��M�6��}
>?�*���d�s��0U��"u�榣c�o��m�qx��H9���Ѡm� <E|��Ap+t
�! c/��W2G8�p����L� 	UOV�����W×C�{ų]�l�喀ව�?n�]��zr�Q�d����S_NEIb���L�Q���,���x*	'�a����kp��V�4R��i,�7�,�IN��������,�H�V�ʿ'e�n�kߊ%m�^�h~5�P�_8OS�,������N�(g�������b7��Lx������e.gA	t
/��6���c8�y�Fb�*;�eq%�	?���r���Հ���n��捵�� AU����1[<�!q��ڔ��Q�xU/�B�4y�lV���߭e�W��$_]ILSoXM��!�x!�6�a]�ǒx:������Zۍ������*.��8��8άB�KA��>�Ht�{L��P�ߔ@���p�,8\h\3�1z@c� �!��ܢV��̠`oU�!9��A$��wky��ě>���w��k��R��	-tp��JU)�c�����k���y��÷w����s=6�}3L-t~8�B��yj,Y���y��ٍ �^H���Z��=KrD\��Iw�������w��1G�<X���J%'��(E�Ӛ��vW�]���u��EK�O�)mT�Z���Ñе`h���ړK1P�/�x��6a��gG�%α�*�E\]<�~�ɦ�r\'�L�ɼ.�\G�[1Y��Dȝ�"�w�-���?��W�L�K�LWP����*���`�MiNy��$)p+A�%�E�H�� Ic�pY��H�qu��b��M���8}޴��t%1���3��164B-8D 4����l��z�'�T�.Ŏ�BA��b�����}!AJE��v�Դ�>s��J۪|��3�a^9{��|����Udp�zS�b[�u]iY��'q�E�Bh������u1��k��y�m�Tゑ���Jrjf(�[�Q���C��[W��ي��(����D	��3�$[��H8�� �<bx����ݵ��rr��d�O��y��8�q�r��VNA����$��UЙc�TA�D#��fkJ4���Oc't^"��z
E�zp��q�iA�^0�29P4��.NEi� '�B�ʓ����w��Qs�+;8���'/D�' ����k������(�չ*J�����|,���D��&(dSj}�(�}�l����~="�%���,Θ�$�ݷ`U7��
����c�.�	O�{���-�O�B��<����[��#��U�L�s�����q�Wb�}��w�ӈ����ӧ���4v�z�~�N�knnsI��:�3����@����$��+���fR�hα�̱�Ў�5��d&$_<eG �o{ං�ü�����ɼ"��k;ٯv�ڹ<���K��	�/TM��O['��X�	�ʹB͚pi�������m]؎Y g�ߟĴT�d{ƃ[cW�@8���e��q(՝�H����G@Xy��S�W����(�������mc�-q�ΰ�h��),'�&O�J��ٿV�+�U�@t��Ѕ�K����c���l TUg�ښL/S�U�H嘡����˺��_������g�y�A[in�~	�@�롡�nE��i[�<a�qo��a#ҳb�������R4Z�Lw�8����b݈"��G�v��D��3�I:�{'�3�1iG�C�����gGr�g�h<Ȃ��s'�u���y���� [��3��������T!��`��.�'�ɯ�Ǯ�y�*�\� �� ���{���ӱ���"W*hU!4]����Oaڳ-��>������+fJ3�jC�~�kQ'z����H�)҅���o<�TuD4��E��Q�\��>[Ħ����f}T��J5c�e�#����������!��?C��������0C�z���B5w�AG��?	��oF�7I�}��W�)WSQ6^5{��'14#+�����AkС�!���f���m��,���0��C�-����^���������j�Q�F
�;�R���k0�i��.�=�����<d{���,;�������VG8��]�0FE^G�A{�oy���@�!�ɛ-]������$�۩B�>��W�A@(���&t_����;T��tIZ#A� ���� ��(�N��^p [XZ~�{�"r��w���!�e� ۧ�]K�(e��g���� �
��\���]��eH�t���'�s�*��)�s�W �E��I�q@�B��["U�o֪�F��f)��D��UλwRaXŘ�������v �p�/�n �߃۵���1:�Ϙ����v}��s@�Ii���R֣b��	���'� Av2�����ٵ&�~�g7�2�P���ko�.����fP��u���O���-C]!-D�V����,I���[*�G�����Vd��Իgy��l���ld��7ו'�mp�$�b�R`��XGn�o��ԄWt�/؉쁉ݱ6����3f�����=���q��Ou�t�&��u���w����HI.tF��{�W���i�uk��O�<�Z�@ ��h�^s�کӄ�5����Z+��Bsr�|�4ˡf�"B��F�%w����f�38Q�H�p�|{�\�q���i�Y����I�	f"X���0��=�Z$ Μ��{i��	&�DL2Q>��Dxe������G?҆�d���ʌ�o�B�)�O�2����05�YV-Ml-��MS���������a��H���}37���?(?�9�NT��X�H�<����XVMk,(�u�E�pCVZ�*��ƸR4!����Rɰ�nƮZ�ӊ�����F]ҋ��k6hIg�7�ʡ��4@�#o됳��\���� ��
���N�^XS���;_��'e�d$Z�
����,�P ��J�8�>��;*>�w��M6*�� ��X�Z�322��5?�/nP=E<Zۗ�3l�yؠp<�����٣��Y�iC�̲��N�q$4�4�%"2
PH<�E�Q�TM�>��zG�Tg��Ye�#���Y5<�U�)F[i�̡P�}yp�YԐ���L]W|��.J��}�0�\�t�a��n
�jgOo�B�F�.��я}���q0��t��`����x���b.?��C��;��"��_Z���N��_gU:�ֳ
���^6��j7ieM��|u�^x��)�O��r�8 7�����&$v���Uu�t�w|��_&"��T4M`��Bu~�k�ט2׺��;-h2�c��~�eky'���L�M4��A?#<�O�;@��j�a%ׯ�%LSh��j�:���M>]���7�<c�V���"�5bC�3Jgm"��P���R��pڬIܲ5qX�ҞC;�[��CٴmR;��3� �b��[�p���[s���eO��v��\�z s`:'�r�y� �e�܋��'�sRI��]c��ryW�{7�-�w=����_��'H�ob͆A�6_8�tT���d��ºbi��J-���C�^WӘ�0���N��-���#'>�F�k�	��#��~��#�d�D�$�h=�Z�X�3�W�V�'㊥f��pK�T��ϩ=Mg����,p���"�;^��#��p��<�֭注��Lב�T�n\&����Hh_��e�\�5lb�
=!�F�S����q�Zt\ri���x� I딓-��Ի����KHОc[��jptBE��%�E�8$m6KMq1��"x�C�Q�u&�0���S��(�K��פ��Hft狮,b�s��!Ud�w�$�r3���/���J TG�(��^6g+�7���d� ��L~P[�vc49�%�I��ƻ���{͙�i�u�I�Ht l�A&���
	�#���h��i��4��[���	"�Ȩ��n'5}lTZ#)�Z:����V�ev"������uX���C}Te���;�5q������c��ļoɗK�D�͂�z� 4%.�.�1p�;++O��#��G%�B�)J�&���F��r���6�~�D�'"�@2�&�ȩ���թ��jw�=���e��h����um�/�^Z�=��E�#l1j�7���'��������F�¢�l��j,.��h��TC#0f��{�n�'����x����oTv�3��Yd��]%X>&����ܰ
�jO8>R'��y�.�g��E4ݱ]���Q�xW\ZsXΉU���Ӹ�v^��e��g����y���!U�yk�ͽ���u�h�@�FOl6 P�mxĻsؘ����j�QDi��D*��R���x2 ����"�N� �>u� ���o�|w��b�f/�0I��*����ոf�kb�ŷ�$,�_�h2���K�B^<�[���̲���Wn5�a���Nsy'z?>$GG<��`C�)�I���k�0)�R�RXo�u^.�S���u����HJ�|���f��WC(���l?�����q���-�b8��%˷Zt��_�>�qD�V��f Q�.��{vM��,���Te~*�������n�XhVf�s*(��'��?�%��%�s�NWH��$P�I�]�M�]��c�R��3�G�ܔDm?0��f�W0��L��z1�8�Ӂ��_Ɉ�Ծ�iO�VM�7ģkn}Z�Q4���H�W���7��[n���h��h��&AZmY��mQ{O�(ψ2���_r�|S+c��Z!B�h�Ӵ��jH�$�^8�F=�<���DY��ع�����,]p�����9��Y$}�J|�WY�9�b��T4�n� �: ��������
AG�S�v�W:�ߎ4�)~k��D!��V�o�R4g�I���z��4�]�����qĒ-_���0!;�h*F��g6�G�����~�p�.��|�f	[���D��O0�K_Y��q�"�K>���IM����$ct��E�P-#��5��P�q#A��ȝ;�x�HIw#*+�&
ȬG�׸�����P	��b���q��u1��O��E��C7�hD)o��Vނ9Y3k��#�`�y�y���V��Y��K=�~c���q�y��U�!�'�o�RZ�W1|�8�?8<>ّ�:`��	���P㩈�qe��wu*�7լ$���F<�AH�|�[���zz=J
������1X�j#+ܗķ�Z��M��쉘�Հ�b���Պ����mxY���,��I\����5�Vs�Ĕm;��.mgF+r��ԃB�%J��e����I��X.T���F�-w��"&�:�HOX�������C�s��kZ�X���e�������y�wE&�<=׬T�l��=�XyĘ��՚����re�)em��^�rŔ��@X��Kf�D�w�����.G� ���1�t�5�+!�?$�o`��e�1yH���:��ׯ8Ӆ%�a�����EZ7<���0"l�Ϥw�K��2^�/?Hm���ѳ%]�~%���c�ˮю�Ʋ�c_�ž%��z�]�?��Z��27�Eӎ���N(;&N��!ɋ0�n�ц�m�+��:��לE7�Q�fws�x}��n�f��j�)𢡊`g�L���Ƈ�j�+����)���~��� Β0��DMFsp ���T��E��B2��`��e�����+�bZ�b)k���հ6�*��_�����(�h�Dy�C ;d�����z*=`["o�8��Ka��~�-�ڈ��T��F�$���Jqe�6��A������f�K�N�����ɝ��+������-��$��&1�n���f�� :���~�,�Y��?�`���G���������"�;S�,�!xʄ����!n5DI?�	��1� U��q�<t�D����J�V�j�(�T��O��d�Z���3�6Z��KX���:�qb��C��8�U��D���=�ſWt@�� yD����j<G��e�y���a�$�5����n ���D��Qy@"����Cu���K�>���k��J!I:c]D| �Tdy�
|<��YNNq�q_�?���3���j����鬽���]���H��_��o�-��$���N¤���e� �҈sw����Ơ�e7i�j�B�=���b��~^�p���$��ώ�gɉ�܆Ykqn��Ĉ����v�f�ңxԩyݶ�ۢ����MFMt�_���]|��ag�<_ Y}�ؘZ��b� 	��b��>�8<��I���6���F;���~y�G_s���Z#]���
��}%m���/v�1lB�I�.���;{+�@Q2�Qхy�^<F$,�c>�T�J�@F�,ψ"݁�1Y��`;.}�0���� HghK��:;���8���^g{V7�[�gfJ�,�{O���f��ҩ\X+��C����m���8d{�Y_ZH�Mu��5�'�^'���L�!�\b�Vb���	�et��SH?�s�3A����L�-�a��~�&)�a�g* 8-����2UO�m�z�Q�62OLI�"��8�@�q���ew^��B̠��6`'$��kx�Ņ�W'�>�Ćy�=o�����pu����6D��.U�:�xu�_�d�@y��fF�Đwr��������A�=1��v���G�3ʾ��RA�ɓ�.6�UGIx��TGl�b��n��j�^�LQ�ҡg�������o���җ=`��3����YE��u���Z����
|��g ��m�JY�%
4�SOfx��6JH&>�\Z��@A���<g"3�� O������W�YHc�E@�ʨ݌�����e�=�N�fyO��V��1�md-��&���e:���fy��mj?,n�0��?̄T��k+.zM�3)mS�1��'g�Hg;ւB!h`됗�,z�<�ϲl]q��An1ʧ���eZ�a����>�p�G�[ϱpBtN��
G��O�|��0�+�,�xMp�	a�w�3�m>��%�h[��&LO��[��5
fQ ������iI�-Ҟ�G������ڄD�������'W#�:Z]QR�4z��1��6���y0J�qN�u%�{}�Va�x7�8������86���=�m�|*u����c���_57��}�rd��/����S�@J$����$��Lq=_��o�X�E�o"d,̮m�ۨ��RiZx�1!��d$Q�e�,�_r<��qD'��]<���y�K�G���W����Yt] �y�Ӡ!3~�h����jR�3~T��a<����OJ<�X\�f~�,�(���O���f�u#�m�E���*/��qZ#c���(ҍz�1*ˤ�w������?c��ư�GA����mnXMEdV�(�yxͰ�7�I�ƍd���|'�W��)o�޹������5^��җtk5���Wy w�]מ6A!v-�v}yb.D�s� �m���v�c��2 +�T-�3rƐ�Z �r�Y��m�"��B|��h�[B�&�����3;�b�PϷ��s����X<�S�����4�렐���Ғ��/���;��0�Z��5#l�^�ʋ#�Bm��]�o���I3�I�c���]����I����hh���"�Z]ϋ d," �Ԥ{�Q�� wK�=]����R'�E�I$�x�X��	H��V���H
��F��~��'\��<��&λGz������|@p�o4�2����UrS��K�?�v���ǃ}_����a�`
h^��a�&)'x �T�����3\��H��B�[��gܩ��O�o1��\��G䗉9h	����?V�"&�*�I���7�r��3���I� �rO�)Җ��X+a:� ���b�"��ޅ�1q�5��߂S���ٱI[x��4C���c�hv�EN������{���E�,���:��r�b�Rt�hA���$洎�^���'f�B
��>�'�35�Ԣ�^&e�CH4@;�� �r�ڠ�-�I�]�X��F��IJ(�� ��dm!v��8_ ,���f3�i���A����}gX{�:șWpT����m����o@��mG>'i���@^ׄ-Qm9�`�Z
ka�^$����5wʮ	��9�j�P�M���Ћ}Z�Ӕ]�8�&e�G���;@�F;!(1�?�ߕpy��N�^��]�D��̐�ZP\�aBYB����֥�F�j{�����Z�ί�被Y��󽯫3��o���uȡ��.��G�h�
K�ؾ�T���i&����k}�+�e�"�y�A��4oS��;s跆�,��C�_��
䷾K{��Z���*�VR�ߌx /��vk�R=5Ff��3�

)��\s�T��e	,I��fg�)�'�Qb/D�����1�J����J�$��z�h�>��h;1������3'ך��
�la.f�����x$&�T�/9��bI]>�җ0\x�)���vX��1�z$aS��E���^N��kR��&z�_��;7^����~%�%mK���CA6���B�,��4U��Ձ�v+�E))6nxс��N�C"�1��r��"6t�%A!q,�d.���e�}i!P����s?n�q"��,E�)�E��� �Y~��Dp+�3͍L����ųӤ�A��eS��N���B&�;K��|bW�����=~F�m�1I�lj���������bg����8��-���MO�G0|�A�m|�:h�0
�O�al�D�0�@��|Zv/��#����mG ����k�p�ҋ��U�(Kb��l����x�˸����:v
�裮"�0�����4h�m���7��ޝ��5	� �W����ʩr�:�N �K�%��٣5� u�u�Rd�t���`�QL������uSi�'���j�	�#y�۝�k���K�����wE��#�-��@��1VS�}�,Zx�ĩ��.
�V�a�/!U�!-����ض}��8YF|ṋ>އ,�S֢���{ɺV^���c�g���=*D.߉��`��G������0ЗϘ�ր C<���Y�5����A��lI�
����U5���JLz�����P?j�+*L��zC��+�{_	_�p %.u�\���@W����(˵]N`��L�4�������95��t�<ַ״e���k(l�|/�f<��2.��Mq+PTG�3Sod���Mj���w/}<� A���U���:���i�!0���k���GJ+�[ -�=%B�$�ׁ[�ؼ�׌������(n��w�i3Z5Y��Jܡq�5�z��X����#2�/o���Gc��WnA��f;@�粛��w�J�o�{���}��,C�x)���67%�ƴ�2YB������	����QZ�>xҁ�OWg�}O�J�����~-�Y��� ~4�Mu�0A���|+��j���u��g�C��c�"C��xq�IJ�3�Vp ��k�����}���W|n�w������~�X�*Q�����j����x2C�dخ��.o�n��Dhv�A�_��L����G�־����jM�xy+����~z(�2�r�csT��݌ԯa��d@�������\ ���A�1�WGglط/�$'��,�kS�5`��~�1��`�<�Y���N�k�����W�{|�)�
�J���xBv�6z6��_��ҏ���*ӗ\[�z����}�%���,�6�?�hcng���.����/��L߀��k��7���(}�A]O8� �d��eyA�[�GLI��鑟�&��(Z\>�qV�Bf0z|Ć��L�F��8�R~\}����ch 9��b�	����pa�
�-βb��DN�\aw�`V������ �Vb7|,-�d�������TD��n*t���s��GǇb݂�tp�S��tC0�.���?�#�-�e��3K+,Nf�����ZD���X¢D�o'(R����D��R��q(f^���Z!���5��.���4�_7X�>�Gk7�ӹMiH����n]��E���V�s����B�_�t�/h��Y�-�_	Ltؔ$:_�iR	�����/� }�s\�<�)$\P��8&�,F)|�ݣQ_~cҩ��.Z��(4Q"�І���S����5clRWbvH�xt::?5!��q"�<���;$ͻ�x���a�_���Z�;�� N ��Zm�yرD�ր[`;Ex� ;"h��;B�U^ڻ?I�'n2J��mط?���xKJ[���e�w�#�����[ ��:_a��cA*�TMU��$Q����(�o��Ag���3��u��������_v�I�W\��P�S� c�uy߸e��iQ��r���a�kL�׹?fv�d�����"A��}�]��(V9]�%3�/�)?v�A�߀[_j�}獷��Y뻡�:P���>�`�@��Wp ��P]�5v��󌼟�ͱ��Q;f_�V3]~�a���+�t�"18�ҙ��\{	a�f�JD���Ε��p��̯Usp��q��X�TPX9�=ݳͦ���ǉ[YL���r�vY��T'����5�yλ[������?B�-�T�1�@{jD�N�㒶6�L#z�yb�F�qq���/;�dM��,�k��7�m�G��r��~�J`�B���؜J���f��*-�-�-�����PG�zv�lM@󭟼\�g�<_�k���MQBv�0R��E��76c��4���V�S\��s�lm[S|�{8�k�� �0X;���.��@�\3u
vw_��#�d�+��`�	 ��E�7���{�	���bE/�)�b�$q˻7�{e�p29�	%֕�1uE���w�K��2�<���h��{����o>(�<���ۮT����QY~S҉ܷO�5&?p�0D�<h���o�.���icmAQ�b�5P*�����A:���tP�~x�W_�����	ֆ���l ����:{a�m��z���V����X�����	P5\��h�{��2Lٰ��&i���5@��A�nHO�x U�������fw��]4��[~?Sn�����:�(��3�t)V�1:�DtE{�*c�f�������0�����E��;I�#���Uڅ�7�Ã�-�w1'iO��FJZ�.��B����i������N�&�%!Ow��_�rم��d��隣�-��!%;H�3�Z��kT}^���SB�=��/�aQ�O��U��z�Ae K�{7f
x�7�]C�{PO^L���Wh�[*6.��ߐ�v��mT��Fã�el�ۙ�I�3>�G����+4�v�{Fn/�z2PIށl�����a���'�lyV�ڨ�Y�0�!o�g�{Yq�r�C|�J�ȁ&��V�X�kn�Iso9��n����C����G�����gJn����I�������RI鋝?`�
�b^Q�A��0d?�g��
ū���S�T�i'�]M����������C	��ƪ�b�`��F��;�XSn�gO�~7Ъ{JKy03g@Ƙ�cID���O�@�&�1�X2R���B�)rd�釐�GX$ ,�O��g�`I�-�Y�c�?:O�u�<�z�P�+*��H�v��n��(
?�e$�~Q���OU Z�5��X�y/6�ǖ��	���Gp�},�ċ�+2���"�r��^���I�Ycd�α�����+4�����#��r&�\�5 i
Ep��/����p�E@'V1��-m;�
ԪO.2iT0�Ǽx�\oe���e1B5��0�9H]����X@�xҔ���3�IN��E�R�B{�	�!�F�{��������{�
����?ekȢ<�_pEw��[��������h�Nh��b��af�w��x�~{F����������E�B\�����Ž���i�v/.��1Np����6i?p�;	u��gr�"�gSL
S��^-Y�wfr�6V�,��;�s���hu�d����{̂�j=��g$��s�bsN�u�����Cy���d^�Z�<��,����wj�'@�x (9Ĳň�
�+|`2�K�!��M�#!�� >M&���C�'�����e&a[o�-�ȘP"��4ہ����݃Z|h�(��pa	�jB�
>�n�m3�B�\�� ]CY����t�������8���9��5s���x|���jo�,�G����S�g��P=G��L76�+�eA��87�iX��s��-.zQ\P�����T�&�Y QV�eGe~���Υ�,S"����l:�mv}¾C����-ݾ�(��v+z�C��j��v9�?q���Ӗ����HR�b�𰹦��8��k�H�`O���5��t��=� �N��u �\��&�.�:_�f�-C�E�	d��[A����<�
�'�d�s3 �M����ڀy%�c�)Gv�k������f�֗3+�m��گ�/�jV<"���@�e�,��3�ۏh��?� �,�F����A�1M����f����Q�Q�%w��C��=���ѶX��{/��k�T���Y0{,�(I�� q�/�`�b�C?�'t�b��S̰�=��Ƙ�~�Ŭ��L�7ΎRr�d��}=٦�I�jׯ�,���<|y�J�t�&��+��l����F���~=��,�oO�ҵ7M�5��v��s�Q�*OM�y�@���:P<�^��A��{���P���x)bT-Nݢ�d:���W���f\���ŋ��� �$R�a-|����ڿ�:ta�9�!�=���.���NBq_?G�-I$�R�K�1�X���Jg�;z�L�?�c4���;�o������P�0o�m�I1�so���}�J!�L��Ԋ�!q=��+�
9H������4@e�ۄ���c����(��3b ���R�M��ύ�;G�Ъ��=��c�p����Ev���TX����㉽���Y����u@�/��4�R�Y6\��:�I��#�a�oY X2�`���ۃ��#>�����e�<�����|�nI4�\>Vp\Gf��F�����r]�O!�/&���6ь�FJ���|ƞ��U�0�@'�[����Z�Բ��GAIA�ۓ��kfe�٘����q ,�|����y���q�����CN��{��3��;$�G����{���|E����Mǥ��6Jϱ��,wuq�]�Ⱙ��b�bp�ϳ���%�X�_;q>S~D��LdNQ�
�����T��~��r��t1��20�D&�7{�Y�尭3��d��0�A6[F��5�Vv�^��Ry�r��m�i�7|��ٮ���r������#Ow���\{��F+�A�	ک�m��.x�(w���7t�,�a/�n B�F���_�J�'9���?6f���%���3kz�ÑA�T��	�#���'R�*eo�or� ��ig����=���5q��t�h5��X�ej��2�e���PV���q���]��7M�4Oͭ|���mP:���.w���c����ٹ�>1d���r���ӛ�V�]��k�򝷯pu�G���G��g�=�	�P0:Ә�pkj>1��e���l���s�f�̸��f"�K��T	m�;���hV��r6:5J��椷r{�65N򵘢 ��p�"�M�-ä��	h3S��?�-&���l�:��""�����Bu>�~o+�c�Z�#-.�}��):}=�4�8��L3����ϝ��嘖ҤOVQ��[i`�a`�Z\�QY�A` ���� �����.�.�On ����7��cd�">���f*���_�Z�u��{Q5m�#V����"�?̈����`jkK��r�R��bG~:��/���)�J��6�]H�i�!�;U��|"u�S�׭�[���*S5��@v���'��&KD}�S�&��?r�+���!IK���CS�����T�la��;�s��2��r>�\����<	��v�ye� ���H��g;no��I��jL|
��A��.z*�6�Hn��9鄜b\ ��9`���: `V�?\����Wa�Ogni���q��t7yS����|騰����T��!D_���=����}���]е�L^F����*H��z��8�+�
���� �;ɸqlw�a��`�w6���PG8nc1���Z�xsL����D�h� @9V�v+m�G����J�D\Z��QQ�t�k���;q�RF5J.��q:��8q/8�w�[��F0���n���5f�;B�G8�Fp��.]LS��i��pR�=�h`���1��d�q�vm��.8����x�>�Dt���4��?�t4��?5�Nb�ޢQ�)�D$@e"�I�B���W,o_�Y��7���e��\�S�A���ͭKf�9�R]� v�ր�bQ�����|ޅ|P����C�-͈N��<�Pg�#��94~�iq�3���+v��7{�;�ŏ�z���q��;�h�H}K�Um�c���S�Z)�����{ ��+SK��q�=1����U���Ý��-��騏2�i���w�ٺ�Ir	�ԓEФ:9,C��H'�D�h'��oK�g=��"'�n\�#��i�Q(��@���;z�fo�T$���H�޵ߋ3���ؿ�퉂�uS���e��K��G�J]6Bm/�d�Y�h�Ӣך�LaJ��Q��H�A���h%<����
ʠ�c]���R�A^@�<�`��'��~��	����ea�Ѽ�H�a���8;�ĩ?�O��H&�} V�&L��"�f����H0�w�{,�$�cY<q1��0��"�}w���c����N��Ld1@�%s�̖����������y!�\A9
�%Iᇯ�s�`��YH2�
|�����Ų��b'S�%��?��#J��/f�ǔ�pC(1AXVᛄ�"����؛���ʉ���\챭� ��z��
�=f����<�o_��tX��f��̱
�6S�T_�G����H�C�y~�a�T%N�J�7id�p��_PT`~���?F1�xi˦^�V�d��v�s���#nP�����"ŚhKK�<�n?Ӎ�#�k��;ĵO~�f��~"}�\��1c86��� �	��?�����1��m�m����2J|�!�_JR�ܼ
��K�tg8�<�.챪��[{z�؉�O�ޘ_FN)��hۭ�*EbV�@�T*��\V�g���f�ڲ�M�J�U�9K����!a��.�9�9���ZVy)畵0�����ng��h���p!��]�TG�{� :��n���K�@1�CK4�-�����ٲ��r�A�4?�#<܀����x2���U�sr�������0Q��+jPJ�D��]�ܱ�YE���uȉl�y�)�}�Z_dE:u$Y�7��aݷԣ��E�<�~��w-��f^���C��͛/�MkF&����&��I;�?�wVy���Mr��;�"[K�9). �H
��\-xQ�4TK�g��X���+��#����l�ꟀM�r���G��u~v���<��� "t��˨��Į m�m�'1�����<[ch��FQa���{�� ,��T��� U�>�1"���]#}m�9�wB�-�Q"�##m>�k�"7��<8�R�=���p��<t�'Cw��f��l(�t�68~JOi�L�u�V���o'��H��M�0<k��"����,��&5C�]�ol�A��SL~�F���N��G�d�>�h��q_g1,��MS������E h��ҙv׬>N�p�`���e�(��l�z&I:3���L��8֕�F j���^�l�&P8�Iѻg�W5m���`��H]ʫ`�)(/`�c^y���aPY���>T�4���=1?��m���0B��e�?$�j��ޝξ��Ş����Us���P��_o�X$/��� �xY��=1~� ǑQp�!��20�JC��x�O���'?^�^�z�e�0�ix�x���p�jHzk-^��@�N[���g��!M=�0���'���3"'�Y{�9���\H��ׂ���jX���%� E��g��c�q�o��};�M��8����mxN*z�!��"S�:��wG
��C�йK�ї3�n[��Blw{�!�2c� �y��y'_�YU0��-���xE�a�Fz��L���\���_S*��J��C��{,QS��'6�&w�k~��� 1}�y���.�d�7N_S(j��A�0>�Vΐ��h~$\��9[�0s߷߮�(���fqNn�H���"*Zz�ZNv�NKư��Q�C���[��fC6Y��n�x�N�Е�;%o����0�I64x��������P>�<V\��i�сGf���Q+i�� �J�����sH��Ԧ�r��&��٫��v?�4������8���Xg���W�?&�ޘ*���j���z��z��X���� u��:@!���@�*}���Vv���TD|�i/���=������M\��Z�7"J��-����@+��!f���a��q�0X���omx�;���X�WW�������z��dIP�d3F�z�.O�SQ���N���Ga}X��I�~����E������8uz�I���B�%� � 0ۨsb=2N��簂��c�8|�ʗ1]��_H�
���b�5�w�R@�sKb�N�%�
�׆��5�Ėfh������,O����x�%!p�z�mQ�oͺ���<���
���l�*�C-��-ӝ]�Fg�Jaa�v!g��<��)'��H�Iv*U6�E��ݽ/�~̆�&��p��ؔ�ż]#�Y���-��򰐏 /�4�RSh�a����^+�p,�q1�O�.3�Nث���h�`ʗc-�Mq��R�5�js�%]̀{NŪ/^ؾ-��e�+p�m�a�R�e��X&5c�I�'Oi#U�[�I|E|2�׺���NL.�����|Lv����r�́�*m��BS��.텄<:�nu#e�I ��Ag}NAJ���2 k�nv<��aCW(㨃�?�H|�5"��p�>��'�>)&����|�������������ѺK�R?1Oc��8j���zn��	"���ƅNG�T]_�E��k������b�d��Tp�������>0��}�h���A�;1�ӴD��|��E?�K�d�?8���c���P�	8�p½d�a�r���<���[޳��w�\^wK5萊�L��z�UA�\i�*��^Q_o[�
�/��8�R<7�$o,7p�'"�bݺP�S̨�A(}����\e�"��ׁ��4���0���I�IU"��<7�K~T&����!V��x�z�xa�4S�Tj)2��I>E�K��e�[����4h�g���u��l���V۰)V�t��U�j# �[���v�29�g�dN8u+8�"�}�+�"���Ǩ?����ߺgX\�:7n#f�r�j��y(�VxAj�敆�0kRk�$��"�75w�o�D�ɢ�Oi��Y��]=�Ԫ$*�G���I�(ٌ0��tPF	����)1�0sQB��w������7L�|��J�I�{���6⽙�(��x��̇��8,YgP�n�G-�l�A��~�o}�J�`��=tM�.���X��+�@ZP_P�̓-��&Z��3�Ǧ�F�@��\�����D5[d�?�Q����;^y��KzD�v�A����Ț�_�^tRm��IJ��JQ���P�+1���S9	���cR	�T���	�n����fȐ4��Yg+2��"�v��{�a�X�,�K��x���w��eD��Ѹ�NC(G߷+�O�uaN����z�S���B�Έ��^�@i:�U�	��m]�8���qh/jg�s��Wz��ړ�k��n��8:�����z�`.�\C�[1ԁ:'PN���U東4��ݳ\�4:����03
{���4�Ej҈Yʏz<�f���^7�zx�f�GlX�M1��Cϟ�,!c��<���u7z~{e�"_����O�ɱ�O`�-i�
�m���xU%� �����K;s��L�+�E��
s�R���R���/5�����X��(o?՘}�Fw())CQB��+�$���b�m!A������+��z��_��*���`��	Y�#l�r�{!��c@jdK2�VcE	�7$ǚ�5a*	��C�1P1Q�XЦ�.+��L^���oft!'�=�[��!��U�zt�F���c�e���R�ycp�a߫tՐ�Ь)%PKF!$��/�ʢ@!9�<�Fԃ[���hA�nW�r|��i$>�}N��j@&�8��-���vӝ��kA�z<c�xU�w��A�4��� �����T4`ÿ��­U)�T�,�Y���]~ˆ�em�0�����%5�@��Eܾ�9+7�Q6q�!����6�PA�[��o.9�D�]�uDA�k
ke�O�֏c,��?���q�Q��dS�Fw[��G*u�o\/۾�77�*8Ui���F�9=���4J�m�������Ɇ�8c�?v<7������R��^Nf�v|(�m��"�Vb����ɀ�����A*�>#�J��aX��Wgt��A/o$�/�#��5w���N�֏��d���-���lԌ��I��Y�+�X�%C�YhS�:� ��2���+:���ڲK��s{6�.�-S�_��ڽLD�8��nݑ"�ƙ3C8l�D�,�B_{��&�o��Qm���I�����U�f�\j����:�Q�W�l�f�Nq���o$^M��+����n��(:��pڹ.���N���?@]�D�I�0��+ބ��,�d1F}�:-��BY�.�2�TmA�r2�)[6�^`���� ̱,�rUo��k��h����ʗɀ�13�I��!���	���(�g1�UU�|W6�ռfK>�H�u�}W�l�\�k��6PW;�|$���O?�U�ض	x���^�p~��ո�\�˻���Mql��~��+�*\F�!�+�
M��N�4��qz�x�yƓ>ط��#��m��S�U�l�k`[H�Ev�M��xG����R�/�W�_
Tj1�������BI��˗�d�-�������}(j��W�fݾ_�A�櫄�,-ۚn:.Q�V��s5?D��d���ˌ\'���1�L�g���>y�3�'����� �ʚg�cP�J�C��g6W������0������V!���vͰg ���h*kd$���aZLp��I�]�x��>�4��R�$��w-ĩ^����v�X;}�lX�bbkK�	`h�=��?��W8�r����3-�w�s��A�U=�y�^PP|��֩���dLX��D��Ω���E������ ��n$\��XS�x�H�6�n��Z��VG"�0�=xMы�wg��y���R����CK(PU������(����`�95�.*�-/�P����t�ݍ�8���EX� ��|Y>O4Y37?��Q��_�V�xY���&`X%Cc�"�x�a���%�Wr���`��$+�u�R�\3zYHt �,����̇��=P��_�2��\�r�:��l�$#�K�{XRX�����u�H� D��f$	�L�\q!�[B��Z�tr���i"
���鷜��`{�9�O Ezk�6~�A$�Ȱi�����X2�)�����v�BK�� ��	uصZ�yM绪!d,��Ujr�$B��0W��-�q��so�|b���N�����n���e�KnI�$u� �j"�*�

�),+�g��/bD/�A��=
x�l��J�h��������l���E��dC톓�(�̰@�J;�<��}u�F���G~rL�뱻�Yʶ�om���	���~��-�S[�P����BNu�����p��h�p�^}�
�f�Y�oSq�=%�H	�'�K���$+|� .�RQ�f?����~��-�^a��rΉ�����z���_�	������f�\�x��+�).�a&�]u�#�ʋ	�)V!d{}L^ˤD&g���rǰ¸�Һ���ĊI���?L��W� �V9h�#�u����4���������o����JH^K����N�Z�C,��JI0e��fD����;-!����hb+jS��PhEΫP$��g�(X�n,l?���Cҕ�A�b��C�C-<L�&�p<�~���;��
����jF�c��ldU'��Y�Q�Q���b�p���2�œ�^�u�sr�P��{��'��`��J��Ŏ�lV9�ݫkO�#E�u�`�>�)P���Ꞇ@���vw8�Z�kϷ�CV~�$7�i���oަ!5M�᭪�70S[�8�<�����B�E	���c�|���s�I7�E�v��YG�f���`��#���T�y�?$��ж	��S\���+e���ˁ�������׮�5�A����S��ྗ�zN:Iϓ)l��cj�IZv9�;�WM�I�]��&�M�'�(Q���{=QPM|�ܛ��(�����6K��)̕g[Yj2Z��,�k��I�|XL4��6��M\l�=��R�˚��[���^\2:������9�9�Hq�oXfG � dՙ�����NC葛;x-A�Df~�EL-.�ǆ.@3k��eE���2�6%�
ԭ�=D�c�����⦼#:��Nri�G�f�a�3�]��L b���g�<Ჴ7:��5v6S#
|�^���%���J���|�p@ͥw*o��t��bR�M1�
`}S� �9L�@,'�+�|�<�裞\�
O\��UrA�/؜��'����c6�=�o��^������G��@Q������
�;�H9���m�ex�~LRS�t3Qu�Z���R3~�ӜR��ɭ���=��!�@��N��{d��B�WWRaɉ״BX]֨��<���0cY�����Gi�3�5�c�h���-6L	�~YRE���`�oL�6����lE��a��������=��ӏIH����Ȧݔ�5 �x�f��`*S��Yh��{��/ٍ-���6���jmK�}�� ����5N/G������8D��A�@aX�+
C� ]�v�1�4=sFԝ;�gb�~�ġ��r}�^�����7���5�K��«E^��㐰@������tz-�b���M�L�=��"Y��Ep�EP�U����j��B¢		�k@�V�@�K�Ț�r��_�e��Žv�Ԗ�q�ӇĤ��w�Ɩ�oz9��ڥ'Yb�8�9�pc0n���S�iG73Ԁ�Y�\��vAw���#�7&��iڇJ@�s��u7c\.�������Ark�
.�y��w�(gT�Eq�>�5 �R<����3���ͭg$ <NOU�LĒR3��<G�)�mbB��yKr��	b�����	bԣd�^�#��N�%����8�X¾ڠ{�&ꣃ;�0��)4����N5�&�BWm��v��n��?���,���*�آ���}'�	������/�����8��������A=~fe%�[5��Y�ۏv��G���o����aD.��^��N�Y��!�����;'��M�FS��#A�±�#�>e3�V��]na���"�P�]5R����Y���x$�i��yg^��[+g��)�E�� ��ML�7m�gty��U����[c[�t�ȥ!��of��/��N?�w�b��c��������s!Q'B�R��L��-H�H������(���nrya�e8(� �̄rY>��	/���눠 ���a��葊n6ޫt~�L���j593���('�\�>�B�ӯ[2H�CrD�|�R	�o�F��B����R�h�H��V.}�fes�;JV�7�s��S�[�@l��X��"�6�z���J���{6T�1�V��ĈED7��-��7֬�3��=�C�G�f<ُ)j\��QU:����#�:����f��=�����}n8��꣫-|�-��e�3�`pLp�WC������������䇋��B vg�`���A��e�(�h�6�V)�C�O��F�'`A%<�C�l��f���[Y^q��dR1nop���n�)&�Ճ}��]��g'�+���p�H�����g��3�胎$����G�8�2�Ў���h�����E�(u]���Q�)Y�<���NݦU�}�e��'K̮�9��J�[�l&�r�"�S��m��,���s��`0�d�g�I�^���붻f_v���Z�����Hj��|{8J��}5K�x�k���e�V�o�[I����4,4_��ȱ�
.9w��(����F"h�w)�`ejچS"�<J-���ҳ����Y�q����씨o�b��"�i����:�;�tN�Y�^oz)��g�U�THZ
�P�[��'�S�th٩�+.*(�Yq6��+U�ɔ�Dm,�c������/�Yݬ�)u��q0�V��#w?bg/돢�@��>C(^�`�͉i�����7�` M#�f�xWVȦ��kxb
��z�o�y\������i()i����T�v��v��M���ò�YK �I3r{7#�+3%�9���A������2@M��=31ýo��� �*C�A���)��'�*4�L�Tv-�8HN;�����M�00�7X�%��QQ-��19�ȣ��Ӓ�,�G�C�˛!
/��c7~3�@m|!�D�?ZB��8i(��ds��3f%��Y�j�:C)c�L�혴n����^��3[,�y�r�>TM�i���	�
L8�/80���Kދ���g��N=�L2�wxYV�$F9��0��j�+>�����U8t��T��H��?��A	�֬J�&�U����+����mR�8l�b�N�� x[���y���5�k�P
����2�$[u�r�h5���O�\u���j0Ҳ�|!~��Q2P��f���]f�B�1��6c������C%��ZQ|[K���W�*m�@��=����z 4�R�Q��!��uK�,��ACfP��b8
�O�0��=w�裺7$[E;�9����f��v`��S�iR~������!v�ӐZ}���
Zߴ����VA8�<5�D�η|�Ql�V�Ib}�X��pb�����lS���Ơ+�8���	k$���,�>�̈����pc��֭��ύ���u9��}t��+&x���pB���ڎ ��m��g��@�m��c��0��:4[��ٕ=�KB�U#��E��!v�d�"�*6�����´�Ġ*bV|K�H2{P$<�6&<��Lb'MG?-K�1|
����IU�����'Y�8�7�Y"]��q���a����r�b&⋒��Pȓ+٨�	Z���#9�����Gjܳ��Y�퇩 �L,7ē-���>9��ң䏔�{��;��r%T�,;�d*�[���陊_	,}H^�J��?۰q2���'�v�N��nBb,�%\��g�d��3���x�h���b��\�f�+���� ��~D֕i�Ș=�D�>�:�+�d ��A�Lk�]o�iÏ����O���2]r*2���H<'�g�d�<�%�zSa𪩯8Y��i�r|C��Bto�Ť�5r���.F�|S��A�C�t�ʵ4K��^�/�s�|�H|���#.=���dC�M�jO(�|=��K��U�{C�mE�$��������c����⿷�f{�C99��T�.���Y4�Y@�l"f��bض0���P�Kd�䞝B����?��Ӑ*"�xA��D*��8n��(OF�]IDr,IW�;x?$��C. ��FĎ4)���XU_��m��C�����?|�n�wk @�y�N���xc󨣤$C�Y�i;�>�b��r9�g_4\2��ʼ%�t;&.b��\˾���*=���	���MةL�j�ߑ"�,[���/�l�j�~��vk\�'���)^嗲����t�>��U$+(1�[Ɩ�6sC=���<�)��~�-���qJ�~��``��lV���\h_q��CyQ5�ԓ��)��x��D�R��0?s�,�v����H����H$���������_��Akja2l�C5�4*J��)�2_�k`>��)ʞ����~�V��[Ia�xr����+˕s�� ��5T��}!2�t��0-�q�>�.z�����Qs�-Lfۧ��o�Vyk9a*S⹷��@u��q����P�կ]H/�W����Y�����3�
ܙ���i�m���cI�y	�S��������:�p� ��O6�*9̥B���$��\S�u��՝����;R��&9$�
N�]�R��2е`�u���B�&F�V��t��{�<o�u�����*��v8��7B�����{�Ͽh��`=�@�����817Xb�*�[/'�I|�R�n	�x&����*?�$�7BO�������zI}�|(�;���+ ���\�� S��)��Ն��q`wty�\ܽ���(cXW����@�u�>p<�ޘ��Kg�ts/y����ʪ�nގ�1x�2~l0�0��🊍�V��/Z#S���[a���ֵz�q�X��F�mV�B��"�~%`�RL�OϐZ$:(�X)}m+c���I�P�[�#Ѳ����������W��%��Ɛ�X�J&��}�-�P�H�f:^�<����܃t@��ԥ�+�����*Uۃ0��t���$���;y̭��������{��{y�"�=�)Ԥf`��XHn�ڶ�c} ��k�㴢J<�w���M]^Q���ܲ(ɦ�$�~�e��˨��f�1i,X�-��f� ��j�."�d!M��m��PՃ�ӹ���
y��u��h�[#�׺�o�"��{E�_a�bu�e:�?�=9�s����|�S�c���	���+�?=3�ZS��4qL8r�͖Q�܁�ߢ.C��k�-�FD��Z���&�|m�:Z��������4l���S�3��ä8z��ӹ�?����,A�*�h
�n!�*��
Xյ��	V)bk�jN �>m�7�s��S��3�&aWjv�Mtf)yO�t�6;)K�SL)�p"#��zE���9E-�19�DA�b韺Kkp*	W�&]].f��34f4fXt>�W��Gz�����_)yTPrߒRY
�.9�y��O�m�MEl�ίq������d��g�᜗s��5+���m��!���i]�{��=%o�S:��lRm������N���$%�g��$0s:2�#l�r�A���)~������h}�<��K�i�c/*U K���g
T��σО�M��-�!�-]|1T�wUţ�Y*�Ec��E20,��H��1,!)�݉0�zy&�=�X�@�`T��.E2&��ϹдS�PC��T�JY��i���u��p�m���TKh��R�&�q& ,�׳�'S�ƶ���d�閘U՘�gB-O(s@��I\d􌑖�-�6.�l4:�x*�0t^��2�^��ی�Z9C)ۍ�;� `5�?���>�e�7'ݲܾ����w�c���K��������)�qJI�/��d=�)%*d�1 ���_�}B/#H���IG�n�����:��'��Rg}	P�ܧ�
��I�`ܰ2��u��u���2W��ɼ D$q5,��1���١��g�.	�OT�'N�rz��'��d)�I�'�){ɥ��m���$.��h��+�-���9�)��ŮXh+�dt���(Y��j}���{j��Ǽ�]A�X����g�U�r�`Px	�-b�בJ�1ړ_R����p�g�\�<���fa��h���;`$�:�r gJx����k�Ԙ|� �a�#�6Qc��+��"�S9}�c|C���q����I:��z��ؾl�JI�C��i�
��&!�OI��)\�S��g̳���>U��&�c�m�|���d�۬Q��)�c��#d+���J]�!���2�6r��o��;�Җ ���2�,Kg*g��z�L�D�l#��xDY�F;,�\tDN~���儝~� ĕ�O-M��m}db�%��9^���b7~���$���U�z����1�ߋC�'+�ŋ'ӺxGl�0�q���d�x�N.Ğ��K��907�ʎu��SU�~���Im,V|�';���W֪�n��S�*�lM��	�bU�;��6���&���/qد�[X\�3��p�u���:E�ϊ�P��*��.�j�cx�b��ѝ?S4j'�l�E?�z$�A�4~�^��w�@)����uY�8�`�!`軕��\� wȐl,#���t�.�̵ظ&�y�6�A�Z�Ѿ�_ď�^[1t�N���}�};z�^�M�oMC�t2K���ZKnuH}�4��,��+	���2�){�Rf��2nyXӴ��u�k)�y��h�T�������Ç~p�ݶ �맿5�4J5�@��#�	�P�pf���0�m�?�����R�?���s���)����mP9bn&�+�"�
����{�kd�{�� �Ik>cX>�p�(��ծH|XX��R�P$�E�~��Lғ���k�#��R���[�щ�(Y�,��D���I��Di@I�j�n�7e�5G��9��C�s��T�Fǋ>9<k��Q�d�2`.��v�`:��Tjo�������s/�y>@iL�`�\?��2�8g��@�=�M��8��yc�hlz�uȣ9#|� (œ�5���\��EB���
\�� Ϫ���<�r�p��æz]�l�or�{ꊳ��Q�~��M����+W�c�+ޕ�����L�H~�N�v�.qN@	 A�\!	���JO_�<����K���J��W�;X�	�hf�Y��`��
q�}Nķ�����i�����7/1�/ϵȞO���zv�S"������Tm��d� 惡E���$Fdrv��,z��歆��=&�h����8���"�F�����6z��lT*w_�U�ϳK�`���7���(9V���Uu�Ē�,�t3d���I���@k��bPS����R������!�z�G�,?{BKyC�?d�U�\�Uל��-��ZM��j�{��ٛw�#�>��|��{�� �wq�B,��KS ����t!����tz���w�g�.�U��>�}D�>�W�+f���{V%;U���h�to�sL�<��iz�Yt��Yt$`8%�*c7��l�J��X�*"pz��f6B~�L��)5'����/�4�������������k�0g� ٶ�j�Xw��V�֩�E�&h�^�Z�8K�TC��oD�����Z	]�]��}�SF�3� Z����Q�ȷ�S����ᴶ{e��G��,��?��������#P���Ϡճ4��?y�к�_������8���2�f�*��C1�PO�u�!' �ɰ8�QB�/ip���ԧ�F�_`27C)�*��@J��R��_7�C��EF�Иc�Vk9Iqj�C��7N`+L�*�!���ˌ���L��9J�y�훥��P�};"2�9]��ȹ��d�3HjB�
�T�1�9�t�O���-�k�����R�*�'v�:i�l*� b���΁��� ��|�)�:ˣg���:�+��n�7��[��n������%G�b[$����}���.<�U����}�hQ�'-�'⮘���YJ9��}����	4dᙶ���VZ��B��+K߱�q��>��|�4v�Mk'P�"�0�Q��@U�!iw.�p�<CC,*�h�"(6�#
�|�(�fsS��[�d��c��z%����B�ff�)�Mԋ�٧���`{݆��1hS�3³<	I�Y�M����ki�+�]�1f%Kg����
*��I���\ʃ{���Hi�w.&��͂+x��ǯ��7P���5�����+G���O����F���)^̮�,
�( �q	1�f��'C+Jٰ���.q�>	� ]��3�te]�ѭ�fTPBb��;+A4µ�h�E�<>ߨ^^�#�y�a��=P��y ]"��.�R���㠢���e}��5�k������$��+o�W�'~5�mO= <���ޥ N8�\gq/B����Ȓ���|5��ST���
��׀q��Q|W}g�j��yC�ڜ��
V�����[~�qZ;�#F�y��c�bR�=�f
�D��BP�=��߹W�`�(b�����l�4u�#s4O���������m�2$��nz���x�̆�����%�f
�:Cp!��d�ᣕ��r�y|*;1�-�����RXz���#�p�D�#w��;��,Ӳ�uHTN��=�}K�OGt�A���{$���2� �۴�_n7"oz�I՜{d6��2s�Y=ЫG
v`����oD����B3޽������|�VD]�흻��uH.�:�xr{�%�6é�\r���id4���e�k���m҅��Zp$�p0
ȶb]_d��VQO�v
�d6qk����2|װ<t=7��I,�pwA�L�E����z؀��rIfm|�fB��� ��*b¨B5���Z7εJ�
�/�jDQ?�aO ��+F���21ㅜ2C�]��c�0��"S"���Xx�
�u�md��0��*�Y���3p��/^�%��׾"�h��r$d�iɜ����უ���a�gSF�f(�qd`q�{��oGӒ=P�>���.ĉ=�[��B��������?�t�ϣz�ju�6U�6�;^���6jd�@���0Y�=���w�ߐ����J%���u�+ϳ*���3��*'���j%�M�3^��t�a�(��'�/���uƤ�a��Ҙv�"����\��>�+>�� }J4�A�u!R��7��3l�w#x8��	���s� ^<�(�� i�^#���O	l�g
�62�����Б�qL��u广��{��n���O���D�]4&5���\O@&������a�
��;��Z�Qܸ�֪R���7����,�}^+	�#��@���������L����BuFp�c�6�DC��l����ZZ��M��+��b�T��c;� �[�qΠ_�WP#�j�Z�DI�B�jI�T¾���}a-�޿�P��5+%�ҟ��&�����oj}����_�����p��q���qK�t����E�gn��g@�����u���g�f��v��&��CI6�>��I',E�Q��J��IHN�} &W�W"K���Xl�ȉs�j���+�b�	 �:`�8�!��Ќܿ	���j���\��,}G��rd�ے���lUG���!<�*����� p[�-<�!HόU0i�ߏ�p���p%Ϊ7�Jێˣ|��K>6��}���\��A2q���Hx�����n�ME�(E�}W҆���g��3�Z]��ʼ�g�L��ٕN�2Ɲ(Z���w\�f�w�C,,~d��K����|�L(KgB�Wd���^l-6Qs��b��+:G���Ԍ�	���7�0cO ����x�.M=�o�!�F�Rm/?�@�z���I�y��݁%I��L����"��0t(�����N��XS5�gN�ʗ@687���J��Q��r��`�Ý#_��o|��
�G��=�I*Ƚ�`�ŭ��"@=ۛ���P��AB�j���Ivp<Z9<To՘�l���+���q����$:��G�����v�?+/&*�XC5�����q�L��?���<i�j�+?V\:O�cv�S�	@���X�[+�
�^��ݦ���!媂�.N�m����� ��F�4l�j4;�=��B	uִ��Vng���MV��V�@JO`��!����Jc����S�[:�S
���Hx��\��������[*���oxЛ�ΒK��'�k&x����N2y>!���85��奩`���S�G�l�!?���5*����p�%��ՕآM�	����=�l�o#C{V֪��b�@vwaS��B�qW��1�ˀi����R�	�o�E֥����+�ӗ��^�6�x��.fpB�}��x񈶾�+ύ�ԥ����5w�I��ͱ�P�:ci�$�
e�\�*��u����r��X���FC��8�eHA�oc��)c�@GԏQ��/�F��T���6�6��;DW�n#3�S:����8�l����2�c�M���]���h���6X�����d�R��^���� �I>������Q����.���c(Q�g��Rm��'l�p��ZT���5k�� wݱ)d��+��j��� LKb*A�-J�Dr�o�#�(������@C�5Z��,�M��4�!X��J��qփ�ef�)��m����̕X}���!�'���?r`�K���d�O�� ơ�����ZmXև��ɖ�2tE���E�����
|ԛTt���o|��uO*g�6�M���j<��X��.�0�C�i��/��R�F�m^�4sݞ�_�b���CC=���VC�S����p��뗲[��9��ɐʏ�XM�AD��̦>��n!��3�4z��SOډd��ڥݴ\����;���XW�ƃЪ:��g��m�R�N{P�
vA(e��O1�i�k�����#^�y}s��x9�[Ƶ���-%�79w�a�n���]�nȕ�����=5
��~%Y|?9��wǋNޖMc��E��5�d�FI������K���	�^T��@dEj*S�L��5�e1�g��
P�7fL�Y6,��v�uJZ�N�)*h��Պr�+��ϴLZ����c:���;��3�K��uҽ��X7|:�/@�WwQ=h�`�"=��LL���F�u;����oc/���r��`��q��-�)��ȶ����H&}�� �bZ��)ˊ_a,�}��X��mߵ�}�s4�D�����=��Cү��酤koK�j���7p �q '�WW�-Mکq7cſf�h=ai��rI]\����Ӷ�xC�Fy�~�ʡmВ��"J��`��g���և��{�z�t���Tg��	I:�D�Xo������C6�&���&��2�4�<q8
����I��(�q�i����`hi&����͇�F9U��W �} iz�$�'v��/�^��hһٮ�-,�GQ��E�@�L 	�1j�ǰ��;�X"���a���)���B���� 3{fA����<��n����"��r�Թ����*�"6�\>�M�\�Ş�[�.+�U]�΄a�z;�����]ŻR�
������J�h�?hy�@�(D��S"O��%�ЖĊ35,hP+�70���k���Z��E�h�}<��0�1j�l9�D�]:Gv5�IL-d8����q@$�8��������k��������3���3���iV)�3�����qR���� �@W��+�]*q�O�b���Tͨ}9vHT�/Ӊ��ɌQwHLD��Uee�s�$���*�ɟ�r�	�"�뻫�`�$���v`
�E۵X-<�,H��)w��z� x�G�������Km��15F�j�� �Pw��L]��,�������y*����=�h��r�ʧY��7`pG�9َlʚj0�]}��/uk���+�0�H#u��m����nu�s	ۍ�z109�cZ)/�s"�r�J���U}/
�{<��B�1[o���ě̡h6n�d�uQ�%�A�ÿ^ˬ͕o�]�S��G�[�[�����4>�1�D2��û��K�|	��Xn��c�җ��s�L~�?\l֍MuY���]W WT�,QX3uP�7ᄍ�pu`�Q��P��u�I��(������H#$��Q�BKy��sa���F�T��[�ۛUU�X�� ���0���4��y�_��ǥ�a���'H�c�v[^ʽ���X?����I��&d��񈣙	p�F���->M�5�(=����|24I�����>����Yxg���u]�%,V2�Pz�;�㳙E}�Mcd��0�2�k%��c�>�'-��:<-�m�7����~6��^�Fg���C�R�4I�Tю%/��b�(=]��o4�ބ(����~.*���0�y�_�^h�6ݽ�2���_�*yO�ne.W0X�4�h�ft��_N�����o	:R��Fpo�,�Ե�`/�I�r�'�KT~��`��:hڱ�l��uݱ,5��?ǽ�;N��e��^�p]��1v{`~(7[�#y���;�}��F#Qr�C'�"0c������[�ub`&���?"�d9�|�l��7�A�Ȱylm�*���Ʊ��97�n��<$��H0��$��S[ï�7~�\���
��0��.�0�Ik̶�3�t0���FdF?���d��S�Wr��a�_m��?Ô5@O�Y<��Ea9)P��݆��D�CZ ���	������Ʀ�h���9����S�-��'W	����C8cvA��ǧ+���F9mȨM�]�E�(�8��/��ghf��͸�4�)���h�5�}�a&��)�r��c!���8$z�&'%��9NZ�b^6���'�̺+�mQ��¯6��TS���6߲)?��V���~�$I*\K�2�Ԡ�=�]�z�f;�9E�<e[-����A"W��	/��Tj�D�+>���@�������5���;Hٿ�J�ѿ�s��rC�����b1�g�=WO�(+ֹ��T�+�݈�F��"�޶�
�(����x�bdy](P8J�0�?�$M:;��dC�.��9B��&[s���k�d��0�s�/{ku��-�k�(k�3M�)��k)X@��2#G)����gv:~D��m�b�/��)�TN�'x!Q�N�/}�y��v��c��JFJfɨ��Z�o^.$�=o=��u|?�u���b�vؒ(ZS}����I}	4�Ho:"�~A�T�Il��;?jD$�9�u%���B�|l����yA�d2�yO��+<y� O�7�N��g?�zB�����<=P�1�ϙ$(D(m����W|�Q-(+y�Q���@�=��&GHͪ(����������I�B88�XS%��N��=�c,�����|�R,Jx|���H!�g��[@�,�Ţ2�T��	�ʫ<0 o[��Ҋ�<�:�Y^"U6
�V�0�e�>��P��	P>�k��[܄"^��Q�b�R��C���=B �A��+>��݋R�2������P��$YV�/�P��n�il�A�ց3'N�$�̄�ž�3F<s�0':��CrW��+q�1��֘����ܿ���FMIdA��=�K3`.���/�����ع�U:�Դ�ªN�v��<�w�%�#�T*\H�N:�p� �s�Z����}����O�IAW�j}���7�5�m�Ƶ�#i**g�ڲ��Ϭ�$�k�:^��U:��~1��=��=Ջ!7o)����f�t�����>U�6���W"]OJ��N�?Q�VLY.�����-\�s���K��Ns��#�S��H��Smrܮ`6&��b�@�#V�*�ݕ��੶�T��m��,;�0͵Ԛˏ+�q��h�v�޹̙�gJF�HDV��j��PA��'N.�V��KP˞|�#a��6�o_�~_��au�]eo�Le�;d���l֡M<��t�DA���]�rV^���N�s�����_[%H�͑<�!	��i������sg����,D8���h��^�OR��5�9�5�=��O�O�$ ]:樏�p��۷>R1P!P�1I�O���tö�<��>}�A�!���F)~�9G�CW?��YR>ۉ���M������G��5O�V�B ~>���;�;k{V���>�lLǬ
I�������8�	U�2�$΍+�99���t��h��AqK�,�\�I�tP�H I�+�lS���:<�=���uX5�����%a�Gκ^�坍8�x a:N/��5A dj`�H�������,PL{ĐiW5�7m4��[@B��֨q�� �M�[X�>W���v��&�UA9���W���6���6Js�E��CSP��(VQ���fq2�V�	r[�d�����o����\���))+v(vH����菼��;�üE}�u+�8��3#7b�����+/��@�[~ ����9H{0i:�e^�%��i�G� 0�7e>�G�N@�Z��C=�I�1T�˶7:|{g��C�_A
	?�|Q{M-����ƦH��9��j�)�:����r��ɣ�,$P1*�7���WL���@t��u^�'=Jz*U}��eU���|wz;�&�G�=�D�ÐJ�~��]�(��Cu�<� ]��ܯ������V~{���;���G:��b��⚡D2����ꠀ|L�1�U��S�χ����U��L�h��?㲮�Nn��F�Rk
ٝC�L芡MQ�z���(yJ�01�����|���Gs���:@�E�5�7�N�g{ �|y@��Fx{�ql��V��V:��mٿcp�9��t*�X�|S�1u��B���̖���f��������%%ۈl��x�����ؿQ�,��d^Z,���+�����O����;!�u�uA�����ifVd`0��}J���M����
*�kP�dI�epVVW�����E�*-�cvh��'Ub��ϛ��gZ����cYt�'�FW�Y����-�=3%2��ww<���P�w�N,=W��cL*�me�+�<p#��O���a9�
�|��hi�t���'N���Y�c��:�ݽ�t,/��8��^^�C��  ���\$ ���pth���N�AC_�/�[��ٛ�� C��"s��[gR�w/�?�_���Y�t����4���?�&q�%�d��k���;����ͱFk�A���e<E|U�m���;�����5b�L�\�؉��)�d/�Ph�D��$�26�J�Wq�3��*��c&Ⱥ�6~����!��H)κYCBL��o�Q�4S��}��Rު��a���9�tS�z舔Z�8���5KH��^������yP���j#C�~�[��P�p�����1ڑ�Y�2.0L o	��.4ʉ�2(;C��#��Q~�֥䭟7�4�c�T`p'��O�-�֫��s�"��U<��?�?F@Va*�w��6Ǧ�`S0�������2"�����D4Տ��� �4�O��auZ��(�R[�&,�� �`�N�ˎh��3�ὁT��7��ͯp����t�hU �eb��;[��c��v���:�tPz9��
?Ylh�P#ܢ:����g����x�*d�l㞈�� ����݆��^d��G�	�Mb��L�) ��}�=o��92̔����dQW��䋄j�
�5��	����_g���]���y~��^�������c��)��e��0�e�Ż,<�$3t���5��;pʅ$hA���vo�en�a9vj�����AdiG��Qԑ�v���M�9������\{Ӌ�b
st����c����S�}�@���>P[��/�j6c�{Qy�-�݋�����R�MWm!�U���������@���O#��+p�U]�B~^�QSJ��H���{��0�,�]�Tj~Bj�t���[d�Jq�\K�c�����-GIZ�6��n&v��j�ѽ��YY��˚4�zz���8�1����s͟�7���.K�Ʊ��m��fD�_�`B�g������Xӽt;�-k�<!��BX���}�KK�����[�ẉ~�����ݼ�DF�큺�S�C���H�-ޞq)��6��� ���)T4�3�/��\�c�ڝ~A�~�I�6��?��~��p@�;�H�<H70���bǠ����: ���
��zD/�,u��H�B���6c�Â���~Ʌ������M�[�j���_jhx1�C��i6uKj����z���!��e��I�t���Z���7ة�D��b�v���C���i�p�r� y�i�o��n7l��D?ܡ�ə���c�{e�TZ&H�C�~:���A�)N���y��w�>O��?�L�_q5i� m�J?�2��zJ[�[ y]��MD����ە�Io@W
;��Ҝ3�m�7���>�sj���L,
���G��/�Ƒq�\G�٘ 0�N��.��p�N�c�PO� \�����L}�/J�8�'����I��ʃ*��D0����7�nD�Ţ����(Es�)����I9C���o=��A�.غ+��X<S� RK���CmZ��|7"NL(��E��\���T6&��}�Sp%�+ 5ټ� [���ڞƎ�E���T�/?�I�1�� �u��BQ��N�`�4���P���}���tO�^�?n�a\���5?�����@}� 6�@H�{��.g�][�� �/�j�sH8�4N�iC@�̙���{�����ձg�w��6�^#��rDg�����<^v����Q�;�t�C�v��_�"$�V"���>�#�v������T%"UmR�G��U+nNQq�fv+���3���L�s����tV�	�W]A�=:�5A/��umn�K%+�'��x������㷥��J�w�+��$���M0a\�Zr�/�ȃ/ю���}Y�"����h�u"������e���i0 A��2"3:��r��K�K�3ȸ�f��Ѕ����q�'�)��8=>���w*����s8cp��F��Ј�+��/��k���C��lЧb�xq�o�;|�Ь��b[��E_���֢�tN���ɹ��H��l�7�$/gߐ��a������j[��ޜN�}���Boۺ�(HV�͵Bh��v@�tMa0W?����K�1Ƽ�F���nh�D��FZ�,��L��Zk�-�l�%�!I,	�Hv�`a��6�$X#��I-�Ӫ5Ez��8���a���D�M�0���>����z�*1�)<�j:Rk�D,j��|��G�9@���:��|Lb>AEϯ1 R���W�T��r��6�#��4�C�ʺ�%Yk�Fi�e�Q_Ƌ|��<Ց2�]�>P���^��Se ��6�3��Ҧ���:6��;��k��O31F򯝎��xZ��G�6�!u��2zg9&l��	�M� �#�]�P�����);1��^1R�]�2`9�l�L� 1j$�Y�h�l��]�q����9;��I2��R~�`I�%��ǹU��f	m.�!0�WWL��ܽT#'�4��z�k�Fö�kl���3a���?�aJ�<p�wkd�]�(݊j�����(m/V�����g&�	˕\�>��]�H'���O���%Cpw�"�<�/��%�1<3�������bd]\�/*�������W?�PRqA����y��_�XPT�y�(f��]]�&�V^�L��ӷ�
����"��f��%�gY-;�������Iy!���2����D���|��^�����K�n�RPc�7����̡���e �����H/���11���O��)���ϗC���fc?��Q�P�^{���<��JIN�{NG>���C�[@"��{2?��HRN�2V��Ұ������N~���K���OP
���	�(��J��2���+����0���1�`l�����0_Q��s�0e����^�ЩzR�>�7ٍ27��M)!	�N���]��E��0���95yy/���q3�~�����'��/��c�4hY��p����GK<�ۥ�� �Ά-�CȣcX��&n��V���BS6ӳ��O�ߺ���X˥0�����w[U{�(��s*�߲�-C��J�E}U�`��
k#�k 7y�J� �Y:�M��5,�zEJPҶ�9��tP�]��y{E�dd5fޫ��'�g�P[�3>禜}�߹�`��f���%U�G#]�H�4}�*7YR�
BNXYQ���	W>� ��ðpX.!�c�������,DU�(s��8������s;��0����xM1�V��
�Qل�D���,���e��>�\���T}eV����Oer�֗)q�m���,�s{}@ʸ���;���IB3p$��Z͸��?��}�ϸJ��urVI���0���U�m> ����{_���l�%�ݨ�$��X��7V�X��'/�R@���i�͖TǦ��p����cM�o��]=�d��A9�����z�o���xܒ/�I	�ϋ�Mu;�IQ+�ڿ��.���c@�(��U��HZ�6<�9T���CpkI��+é�[���le���
�_���m�3�M�f<�fd�
��O����:�� iյ]N4Aq�ϞI4-&�^~+�.������mO�%�&:����B����*j��{����/����!���%����z��	�3���P�[M��=�I�[�Um�(P�ބ G�5��{���sË#밭�V���%0$uZ�?n��R��������|����&c�K�Z����j�qu�\\�"�`�b���7 �8"�~���u�Ff�.�^��g�^)��\��o�0��l�X�������?DM��Q�����˨/;������5���[�O9Glp�����YT��+���͋��3��չ����/վqǯ������zg�f˿�HJ)rL�L��E��Ư{&Q%��zj_>u�!W"�8���I�>!I8�4
Ip���F�[�\A{�?ԙ��'�'���i!{~H nMq8nL�؉hCU��y��ۮx�|Tj ���L��Ӿ`(}�\�(uDB&g4�j��2�;s���	W���sV�a���^	�/j��:��H�o/�nH�؈`D)���uC��[�s�L1���1({���.tP�9u_��6ή�oS�u��e����L�E������Θm��G�2<��c�>d3:�&�J�KC<�`9A^ZN �J}l�"�C��7r*[^�hԥ�����9]>(!<g_?���o�Ƽ�,X|�4{�x@�k����;�#�*�G���U�IL�]��p�]P)���^��ŷ�����K��}]4�||����r���N�8�(ޖ��v�z�s9���n�lF�ɗ+� [�ڻ.��)S�Iڧ�<�H�W�x���s�i��o(�A-:
R�H��s��)�wT�ڏ-s�Q
 ���a��:i{�h�:!�f|.�a-����(YT~���h�sx�mr�s7ʃq��� G`B�-����4��|�d �u��79�?�*�~��N�����	��A�UOݟ}�4]O������$M\��̛2���� �p|kT��
��&_��3�hX$o<ܝ���f�u@g.�E#��6ej��i�f���\0Y?H@Vom�`��v����:f:U�i�8�4jsa��j���^�#��~%w�t��s�N'��
��*�-�$�
U"��~+Z�,�y��OzQ�b8}�{��6[ջ ��Q�`Yc�Z��=���Q�c�_���z����rB��W�0��ʝ��()4*��h��h_\΀P��.��׃W��^�ȗH߿�]#��P�la�p�������&�5��=U�(��!��t��o3"�A��}�_#$?-�<��ID ס�o����-�� <*�X	VV�#�e�B��`�C��"�uW#�+��`΋��ivX�rG���W,!�P�o���2q���-D�
�j�S�~a�}{q�n{�r�yjY�	�S�����e���A`VFb����y2�klsˉ�(����A��MC������7s�13�{�`�-X�o�8�,>�3�n2T#C�Va$�Q�v�3vQ�=���MC��*��%寙�{�l��r8�b�;��#�q��P���wA�ʦ��'\ݳs	��6zl��GB�V���sK��_FH�n
p"��@�U_�bUf�7��np�����\���V�V]��(�Z3A��En �x!�DZR�%)0d7�1���;4 �\��D��� X>�Pd�};@ 
� �q��a'Dv=���אh�n�;&a�䯓|���=<F��~u	��t�sk���a<l��}����rލ�x���X��W���M�����
��&޼mӥg�2��"DFZ�R�H|�rQ#F%�S�\5�V ��o��^׀��0�!b=�9�Ad:B�&�n@�s��6O��J.�#=z	y)�P�������F��$���8$Mk�# �!��L�	���I�Τ���fi�(��k�K�?˫n+9���@h?����� �]Y�b�������� ��M��2����ha
m������7�$-��S��C�Y�Ju��ajzk?Il�"*{f�?�>҆���tJ{MH��o��!,�f6G�^{��ג[D��Ղá��N~$ݾ<����%��D��=�9�HT�\rb|� \oLCä��(���ZH1�Bn��QM3��:�t���6��=M�)�%�L��\A�4��²$`K͒��L�(H����L!�D�_�U��~�!R�k�M�B���_�I�6�����D�;�ɐ�H���I�<�GF�K%k���)������79s��#M6`��羶��^���5���kXL�?�FGu���?u�	�A�T��z�ҁ{D��M����(�cAIV}�f�����3b��0�/;�a�L܇���E2�၎��{��@�%��t��`����޲��"��{oC=x��=&����豂_�k���r]��T����]�R���q!\Z|��S����ӣ���RW͞�S��S� �d<b��.	�C���r]8:T�]Ne[A�?�ڑ^ל��-���=Vy.��ɇ��&��^�S����j_f7���zF���#;תe��վ:h	�;:���H�"��]�m�f��AB��}����w�
V0�4��Fv�[��q��Դ�f����ime����X��*�p�V�'v�����b\p�_��#?�i�B��3��e��[h�:f��%���~Uof���X9/l��h���~�4RF�q삮_ţq�Q�}΄lLwsgw�[��D&*/O���L3,�[�#71��X�@�Y��Z��b0���V��\�n���N���ݎk	��0&mD�Tm�#<�V��0����	��߄��Ѷ,=���ؐ�S�	�&\�Kesa��an���&5P*[�4sY�K�=��L4��	�����X���t!�?O�-�ek���+>@�]�M��`_Y�E�o���r&B�ʒ.��~�"�x��������vHt�R��km>.(<��3o����t�2(�!�˨�a�5]�.A�������M��1��K�7LAO"�vq��~n�H�N)�s��Y�;��U2i��}$��R�ӂ���yt���胡t���K� *j�3l�Ь���t9��K3g�d^�U��@��֓����-��mh��Ϯ5q��l�L�H B����ER��������������9@ ����f���S��9>zNiPnX�]1����_%n��֔^�o:N\��O�d��-nj����1)P�Xn�XV���T�>��t����-:�r�ؕm����0?��4���-a98�%�[iEve����k����l�w�G$�'��j?�w۶+8���ܕ�����+��ME�l�����Ƈs*��Ó��#�A��>\����i��f+����k����l]{�XP������SǘHS�F���~�l�:�G�r�Q&�y�	D�^�'S/����2%��E2>=�]��]�db`�6�`�{_�"�53^���ͨ�=K��V��E���.�J��c�����1 5Ԯ���*d��b�}5a�fiq�f�z����a@���o>�w|S����D�U�a�I��lS�����"β�^���Cٴn�a��}�v�D�>�SqY���J���l�5��!��Ч���:�I�4հ�J��#v�Ђ]�r-��K�W���S��1�E�#Gc���I�n�J���C�����cf�����@�;9�_�ը�~C��1辔���؁k��a�=Qg�uc�d�۪AR��9�z1��\�nL�.�|1��ǃU[���F����3�I,ʆp�$����R50Y��l�VU�H|'���E�v���DCI��@��{������D�0�!/�e��ԍ�@F�^q�ۍ����yZ���ߐUEshJ������"��ȶS��!��ٞ�*�u@�ep;l˽zϰ���a�����iY�6���2.琀G/��6LZ��=�&\��n�R}��I�������#�E{ד���|��?��'No!_I�)$`L{��Qѳ��=Ei������Op�������ؚ4��L[�|*\J:�!�m鮊5+^�z?��b��I��GE4��^���<����X���� 	��n6�a�V���Ĩ��R�{�FY`G2qy�@�����S����j��Õxz��G��Яv 1�l�d�C��\h6����I�����6�sr�tW�|�ږ�;�9`L����]�'9hɊY�n�K����z�M�Ј�;g-*fH����2W����8���C�B�sw4���2~��6W�����`�(�&�����4�<���Y{ȑh�5�J�#V��j�Jxl��P� F��3����8xT0$����y+����П���:s�f�=8�F�&��h=A	|�:ܵ��ӕ2d��G�U��`���0������^�]��͊KC&��c<��ч3̼>��㜲��ؼupv�)U�������y��B��~,o��*>/�yq`INá�ZiÕ絀�n���ͷ,x���;t�;��fd�ا�@[x�B��WUJ=F�h���sp�Z�=�یX�i?d)?�݆�E�RN�1����5H�ҏW9��*R���t�jao��v�|�����\=��KF���+��zt�f��LO�W�{�OMz^�oj#-���9c�hv��&	��o٩��`�U6�kI�յ���8E��Ô��O.�L�Dh��c�����'����Λq�,m����r��,ȯ��F�D��ͣ��l�S*%V��h�[�-�Le���Sp
���-�<���&z3T�r<�ԩ]�ܩ_��z�H����cA���G١�`&�5�0�HS��u���X弜��|z��>���|<%�S]�"�U��{�K��X��*�N���~D�a5�+v�/�MƏ�y��w?S��S�L4Э�ξp'�	|��Gi�R�dU���ߖ�$. 7	�0l$���^��xa}4�F��h�:V����8����Ci����Y���(�	5�8���m�{b˥x�o~�i;�:�� �x��J����ʬ0cm�}��W�8MPɮ��(2�ʷf�ɔл�����"��QB����_�gO�0L=�X�~1*U�\��>��/����[��4�J�x���O?$�����fT��x�)�y�qB���o3��_F��]l�ü&�u%J�w��GS�����r�J{���r�Mxp��#�������?�4n������O0͜l�"E�8�6��2���������q�E����x^�[�F�A��]:*��>�ͧߘ�4[�r4�5��"��t��#n���#J:j���񍦶��	!���/��
u�p�WFm�'��3��M�:�ظO���@5��U{5���kT{Qi�e�ӝ���h��*�����+ٚG��I��Ju���0��I
� �(����O��
��q?&�J�E0��}]�۔�鈵�Zk=�ŠG\M{�x�4\�}P�����dܽ6�K�o��g@�*�p�%J�q�d�f-Bw�ٝ,��3��޴֨�uX@�25�e2�hK�m���f�~���C�K"�Y���/�^�uw�ܧ�zx�,rl։�,��Y�u�,���>�r���7X_����� �,����5���C�#@��~"���^$��MQ���|��ۡ�y�DE)�	�i����Hݵ�*��N�J慪  �_y���v��%��@�����  (�D��H�~P}P4`;�;��<����F�L�L#�'�T���h�v�0b֏X�*�祭]LP���G�����5>��@�F����C�:�(�*_;����ㄹڷ�R���è�-h?��E�و|��#��@aGv��O
2E�Y�9�ӷ'�����W���R�t���Tn��G��L |@��/��B4�Ve�)�Ac�l5�8�5�$����Y�]��i'��@Ylc|B���4��.�К��h�/?�L�L���R�f�H�����4�K,��bX�8�
g�+Y��Q���:��g���rN|)�o��.���l��:$���e�ؖ�{  귮ԛh��u�cvPz4��� �x;+���D2_��a{�	,�	.w�@ӟífa�q3Y%��&j"��-P�Ϟ�~9b�2J}ݔ_��Tz�u�U~W|�Q�u��}��ɉB��Di�<Ƶ 	"�Ke-;$���LI��,�ܦ�����Q>\����+���`��	������ͮE��U?kn7���S�@?f����\�/�$����o��� ,������8�R���
)dY�޾=��A׺�&g�c�h��"�@_h��1�<q���6. ��v�ck�$_.h:- [MfڏJ����ۋ��|Z�tӨ_=�l0:�N���U����p�F��������QAb��ԘwAaQ*4*o0����۴����,������ߑ�p̼�0���F�!-��XD#ݘ�Z�{��²p����+W	���@y�6.6@�E����k��;����ɠ�W�f��T��ksiܨ�6��nXc蓯��T?$�U�s����v^s[8Xz�fd�`�	�TZ^������}�D��+��,�w�n�R���*���6�ݻ��ZHaf<uR'�mt����}=�q�q��vnQ�@r�aDg�D�%}J����:�;
U�#k�?GH	���5��9_V��摀���\x`�Ə�d��j�"�?-�o���"��5�8���:�ۜ����e\o)̅�ͤ,\�rD2E�Q*Y���|����p�/E�1�W�7M���yy`��K�$�z^�w�T��C�)Rg�Rp�ڶjH����H�<<��Թ�4�$�'���S"�&�q��x�\.��5[���Xb#�]o�����1[3���M�r�N���Cu�i]P��@�:�M�¹��,|�j���-ɡ|Gg��C��᰾�7B�+4[�8�g�`�v�'�2T��Q����v���;�Ů���2U%�'_]��l&�lS��,��eMS�<���]1X�Wt-�1(�(���x��p�m�P!��-��Z�(k�w�Xf��O7�T�`��(�d�PTR��ǺS�$�f�03(|��[�����t<!Gj�x
v�:��.��Q��.��bvn]v�%�Q����QϨ,q3��0Xn���Zbۭ
�JDM�~3�A�%G'q=��:3�Z��MY�\���/��p�m�5(m|jC�����["w���*���^}f]o��F(�f�~�I�t���/5���Jr������QJJS2�8C�˸�%�)���$6�J/����z���qvW��%�^�-�|���� �M�xl�^��Ĩ^C߂���q�:|�ɩ?�*���U"}:������m�X2����G4��Sg���
5 ��VL)Dy(�贋��ꌘ���nXt���/E�w{��5s�RP@P#XY��D�	`�E|�\�/M�L��[8e�7��T"5�͛#�!9������/k�0�k^QOωk�:Mw�{�2^��=�qO��X/@IAU'*���Д'���BC����V�+|�YM  
F�l�m]F�9���/5;�?G�|�)���x(_�|M��*)�eJ��t�����~ �z�B}���ͭq֨�W�GM�s����Rj�m��g�>k�G�Ϲ��O�����堜�#�&*"�|9�Dƃ�O�:�~f)��(���s�1�1��[�~q�~v�͹~��\�+�S��ؖ�r8���K�;�2�*tQ CԳ5�N��R�q�OS���١:]����Bp3I�5U�{)�a~O�+��XJ�|_����\��S8�����#&&)����U�S�?����:��`=h�T$�3�^!������sK���~Np.���&P���Ȧ{�HwO���y�c��r����W���]��=�C�;�]����k\C-��}Gް�f�b�8��E�e#��r4��l��a��ʧFE���{���w�s�P�"Z$N�[ְ��Yil�[5��^-�m�!R�@�2�����`�^~�-%m�vY"����qe+ARTy�]�~�����I���hl�i٘�um��(�k�*^�����%{�g�;Du���a3�ț��kş�a��F�^�${|bt����˅�b��ݻtIsd��r��F�Ʀ�������=���X�~�>R��4��c'w�2r)�N�ܱi�t�sğ���ډxCD9vB�<27����8н���ES��􈊵h��bI�����Zxf6�E���i�=�hY��<]�~<�YD}k;��FGj��ъ����E�=0��:���%�QB^[N6�b�l�T�аr������ˀ̡�-��5|:��.�F�����4��$+��`WK�~�d�Gn��+���g}���O}�lE��	���rL�c6'�<�_�%SU�Gߨ�?@#���|=��6�+X�����y3'�5U&vʤl��i�.�yÉ����9��F����䝽�=��)�d/jb�M> S���	Cl�pb0/��#gja2���Ul�7��a��aq�U���#g-�����Y�nr2��{��L���I�=�_OĊ<W��qi����d=�)Ъ��XKǪ�_T�)��Տ�vI?�/S��,uk뿼C��+���f=��N����"��:$,R���̯-�?bL�Jj+D'�� ����#Y��VI� XHS�1�������B!3�N�DC8g�P�)�$p��YX���ϴ��J�ו������K�1T�^�u'��=z�z���#YN�Z+H��>�`9�F��寞�SM��a�Y\���D�3���f��������r�9�(-��F�DE�4Ek-��Ona���������ɺ�. �s�딞w0R@8�xv�˚c���+�/e*��x�ꧦ��v49e�N|{VQ�B������p��X���xS����mF�&�;������)��K{��5�;�t�<P�R�ا�"�٦���V"��k2�y��Y_�\�ipK<�ROV=w(ӾE��RF2�}��l.���Yյ���Bw?��HG��]�U��4|��LM��aR'�����Eo��+����W��Fgj�ܱ)�,	��/�E�r�qYZǾ)�����tGb-~�*-�6��l<hT��3a�-��g�mJj�Ƚ3[(�4�����¬$�ݯ��)�*u�w�G_@A%�G��F#P[�~^�?�C�����t7� Q1�a���x�9�\]�Yq��Ʃ�&�f0���G<�18�c������|�'�{�MX/͑J���C�Q��E�MO����j8��h4:uP�i*eβES	3�ڦ+�7�l�YM�괽Qi������ェ�v�u��`�_[�M��5�랼��]9��Ü���W�	> �A0�V���i��*Cao�8aB���tME��`�A7}o��6��7�K�P�.�d:�󲃵�T�-��f�=ç'azs��ܪuƯ-����8�̒9)��j*=��8e$������b/�@�b6��~z�Hs�-I��5���F#8�j/ }W
#��=a�姖�����G9�q��|��lYcM��c#%b��0̚�#�>���3�}�4~լO"ZJ�mI�'�r.Ǿ��Uc�I�ڒ�؈��5"��⠎O�I53br��?���RC	g�{�4�O�1��z��ا��M�"G`ۧ��V+G�y��?S�YW�570*�!ƻ�V���j��L�Nr�f���I[��CNlTKy��kz�CiW�O%B���|���ȋ��8�k�M�����<�׎F�Ǵ�C�C\���U�P�K٭^6��a~�j)eI)�,����If��5��x�Q��BV�i����!�<R��{�Tf�a������:�ޟ2��r��TNO����p��Ұ3��C�T_<k8�i���IZ�'>����SRָ���m�<$����!������Wc+��z�X!LX�nx�7-h>W{�5|*Q̝aPA�#3]q)�e��s��^����g�:�B��|sZ�2�Fx�|���ƍ��m���'S�TO�S(Á)W���U�S�5=�0E 6���<^MS�{X��_2u�i:��~?Bb�*�XR3�P�;�+���ķ�E����ӾcMU	/���]`�dI�%<֔��2�H��`'������B�>���	�A�iW�h�.�����(Ѷ��<A��2GL�m�WUOr�7p��~�'�p~˻�d��R����ն�z�a�ݬX�o$ZD�Mc�l�z8Ԉ�g�x��a$�e�\�o{Dz�F.�t/Y�W��qJ`�,>��n95�cL��2�)FRv/��ۿ�Xd6�|$/���w)����"��+Ӟ��(o��dy�����o����uM��T* C����g��(�s���Qi��t�����&Ũ��O�3�ͻ�$��`���~�R:���0�����`z�L�3Ѿ%m���D��H���L�(Po����lN�E��\]N�����6ʸ_�"�F�xʗ±����OB�+��m��A��������}��>�4�`Ժ�x;�ɑ��ӮA,���?�~�j��&<أ���t�����I;u�(�lIWXF\�ӂĤ���T��sAA�
1�02Rg���6j����=�H�oyllu5��t�T~��4G�d l�R�]�J���U7	Z�XZ��k$`X�.�6�5�}m	�/��:��M�����u�Eۍ�Ȑ7���g�������X�ְ?��Q�uK@>;�|7���?ψٝ[��t���BvYC)�vNJ磒I� `1��v�0ל�iC��v������!�q�K{4qGXk�D���c8�,�S4`����RQ�B:����e՛�M$1W2�b$u&��&�
��q�Qr��y��T��:ȶ)ݵ��9�+R�%��wt��U2���#H\yցH�d;
������-�*x�a�5�U��'�3��&G�r7���#���a����\����]a$�r��&����m�w�4�l�vx��fir,tuw�\����F�.��$���/�"�h-M�m��1U����/�P��G'���$
6����}/<�7"$�x ���^a�,Σ1ޙr2��9^��P���f��tR��n���I��k9�mT(�χ]�-�-��������ZE�b�<�K�XROM���x�/�ֈ��:�A� ���ġ���N����H��{��\�2���w����G�|���WN"�����V'\ͷ^�ǌ����0�~5�n�v�|V��j�^�E1��3:i�T.�h�����n>����)[�b�v������p��Yv�a���C��#���$��o�Z#K#K_ݶQ�y�g���l��3!�,$�`	q./&Wn�pfJ�,I91�b>���@8���t��I�����e��!�a�(3�,�xi�'S��k×���r�.�Z��ٕ�����Zi�r!���+�B�KHZ�b�+�8_��R෧���u<E#��@Y�ʗ��ߤ�,U:��n,�WE*�PG/�h�¡�)	��6ez��&��7�C%�7���ߺ1���L]�ޘ��k��w�\�k��Y���o<�y��c�ڨ|�����&7��W���ڲX�K!ˍz��j���v|)�W�j?9�I��^$�����V���k&*���K��q[�~}A�5�����4��9Q{���?��(I�9�F~ֻt�ޞHF�ؚ����IY)��q�c�[< �1w�Rڶ[9�==�����ܑVM��{��n�`a��<���H�Y(��}`�Q�eݿ3|�h���L4q�nE@$3�*��$)Q ��0��\�=��GZ��E-WW�X�0
_"�eR�T6�`��i��g��#$�O�9�'���i�R��Rޅ�i��W���g���I��|�f/s�����sO3��&���l��ģ�ô�Y�3�s*0E2�~������및I�G�=4k�m蓍�F�1ª�G�Y���=d~�'OY@�bnC�C�AK>�R�@�$��� .P�r��c����^Ľ/�%��� ����A�r����`�!�l# k%��}O3��x���pӈy�o��{P��F�����i��� �A��Я�,��ccj΍����a*��k}IzBy	���[-�V&�K4�h8��p�m���f�C�0\k�y��X�d�*��MQ��)��	�Ϲ�'���c��������Ddp�����s�~?�V��$�\�}z'l9��%;MH����D�D��A�h"���P񳡩v��8�c�2:�2#��m���2v^��i2o{�uW^r��<�ʹD��& �/�܃�BX���C�H�i�CB���~�9Ă��#ͨ�'��i���,g2�v�_
zy'l��Hbi��F��ژt�	�t&�����'���{Ua�n���1�����^�D�ޫ�e�^�v2��vf��Iy���B<��b0���0DS��Q�&C���rVL] �R�\�Y}�:�u�~���0���ͫ�R��gvk\I��T���]�+�bTW�y�ž�c�@�g����y���Ɋ����uPx';!U���ʻ���cƗ��������c6�ayr�L��+����1B��F(�sr�&����9�j{-��KhǮ�0(�kD�;��O,u�uw�l^�?��Hn�8��g@K��9D�^�nt�ɥz?-nJ�)���pa>ą�˨@��ór*E&��W�����'���
=GzY,#h�X�e��A�1�j�x��HR�r�J�ɗ�ұ�t��	S&~�*L�<<U�*�ęQ������㻰u߶��{����N�u��������7�����^A�c�-��/��P��D�Άz�2����]�2t{E6В�s�A|3�04��3�7���k�#wg�#=��S��8s�u�d��qF9�XͶ���Ѕ�q�~��γ@�aC�����6q?�w���;˓����ԧ`[�j�����A#b's�oɍ�c	�u�&�=ݚ���Jp�]���R]��	nG���~���xDD�v��Z�t�?�)6TFd������RF�b֝}����'
Jw�٧]�:�?�H����>ׄ�l�Zl���ČK-v��pn��K?d�D"M�����kQ&��Q	f�^�0�l�;�:�؜�w_���b� $���a�.߱�#DP\��+���h#����b�b�
��vf�C����b�b�t����v~|`!m�P�NU�)������#���H~Z՚փӏ$՚��,~��x��b>j��Z��lvY"'6j3ƶ�E�j�Nカ�0��ٷ��B=��T�����2��JNA��0��=)�-����������fH�2�sa���^č��)�zP��j �"�,��96���௃`��u��LDp�Q`�,��꽁	`{T���}`��ZŤ�u��v.j�(��?�c+Qy?�'/���M�{��c����I��u=G�,���6(=�k�[�����1� �h��	���%1�.���R��
I�s�� �X�ê��߀��
�_ݯ �v~�CP�;c}�sq3!��)OKFrj���\1�+q쇒h��c��W@��

�������_#��Q�gL3���?��us8x��KD��ֺ=���a��q��˨���ŝ�y`��k��^�Y���X��%v�*(��]�+C��5�c (�Wcl?��"�d�+/aP���*/�m8�W`�FDC�����k���*���U��b����=��@\�+)J���di�V��˄������DC�w2�X+N^T��Ӿq �v0��A8���c��(Y�],Ђ�P���W��@aE�nQ����%P6ڕ�F"��k�u�P�p�������#���Jau���-���~Ks(}�șVO�^�(t�Y�$I����6��8�Ja�mׇ^#�<q� țRH� ��e�SS�̖涊��B"�|��w?�J��'�8 ��~D�w^6�����[NKQ�y�u��b��S��Vq�*�p������G�V����\Q�>�����7��T͐E-	W ��ok�}���P}wM��ny���;�<#�`>l(����bY��`o�/��b�z� ڪZl�5]@����S��/]��7<��Z��ʌ3�u� ���6C5L�9����D������`+�k�s-y������=[���N�	e�@�������[#o��O��+�)8{��ӒK<���d����#e�-Յ�I�l�"����[wΊ����S	f@F�ntt���/޵��m��}P�tq�Fh��҅kؘ�ų�{
sϨ�i�₆;6�zϸ���:<p��R}�u����f3p�}��2���� �(�3j�-=����6��y�	 8S)f�	��Pg�F���](B����+�9؝�WT�=9W��דo�N�d��9�7B��!�W�FC����1�$�w�M��~`���&?/�_���kUT	����H��]��HQfbMEƾ�ƚ��@�W���e�V�S�ZY���D)d�Z���*/nl����s��Y���<������3���܍��}�{r.�9A��?w��o��N_�����J���W�h�������4K
Ļ6d[6���܄��d����9�ү��r�1��������-����r�DP�,�
������t~�)�x�c |�H�o����^��٫X&a���>}Q�v�/3j����f	/Ea�����i����&ʀ��n�֮��y����n0�]�`�0lS�"�2Z��8u�`�l�UR){��p[�@gUc%Yı�|�Eb!+�*T(縆7�r��d�X�W��F���J�}kԮǺ����E�a�ED]���'�5饯����Ѡ��^�mw>���m��)I���úck=3�@�I@E5ͼ!��#�o�;�"��� �K�'.B��|��{���=_�
�XK@��4<��Q`��eN�1B�¦����]H�dg����Y�E�;��tx�e���G�M�������n˻or�.�1��M���� G���Jxo���2�\t �������d|�BS^�,��Ye�Ð����"����i)&�����x2�l��mL?.��>��Q�}C�'�b����%~緭�D"�d�{�ٱ��fb�� 4g�%��r�U�e��gX:�:��,v����a���/�|�(�G�"��mJ�'Q�h��O;%�5#܈Wܧ���4��ϟ�ϫ����!2���4��Vg�v��߸���j�u�)��H��29��-�9��jt��w#OW9��<-c���b������!�"&�@��}4�(�n�}c�p���?��&$��C���L�#Ks����q���Q�̏�I�1x|�����@U���J��:؝r�['l�đ�|!T�ġK�V �_u�_+�
O��ê3p����/�G��~*���s�_�!{��
���2�9�b#�f{��^q*E�T/4���*��XH#DJX4�]%E8�UUNo�K�/�����/������ SV��ꏲ��fa��B`>-~�]+S�6�e;�������P.��R���W�~��vu�i��(������lM������;�Cr�=�UҰ��Sࡄ�mΛaƞ\p����ȼ΢��#<n�u)5?�Q��:bb�g$T� NA��u��u�OoT����$������pon��&L�r���:����y���o��Ũ 0L�_M��g^Jc4Vz���q1��V7�K�kx��d�9#�c�EGL�3�sd�r�/���kե��.���.�v����0(��5ڝ*`W�dW�0�WqQ/���o�G�̆��W>}I�җ��	�!��sa��hx�]x�����&?.������1��XQ=��R#1Ѧca�G���MQ�O�h-J��u��(����F����$�񬹫ʵ4��ޔ�=�{k3t�7)���0_w��DN���Hq4ٰ��r��"�5�ف��Aֶ� n7r�c��v̈́e�W��{�0%�Ue��sb!��d24lC�q�<��.Ǡ�xC�e�K G�:��n*[zs�I�:� ���o����r=Ӄ��Cۂ�Y��QI�s`ߔ��:]�.��� e:����yq�h�J�u{f��Qc��gP�z٦ՙ/�ʂ���pXqx�u�5��kۙ�O7UɎz�|�_�/t��n��BO�g�:P�ƛ�Ŋ�_>�Dd���6�e�5�Ѡl�3vJB�d�ǽ��A|������ꫠb��� +
��H�a��3��'��'��~��{���A�R��~O��y��
ד���XW��˩4$�	�(>Vn�(t��2C_a�Eg*���� ��`�ܤ@{��',jR�N��nbz(X���+Q����v�5ھ�W�7t��N�s�#����j$��W�r��Z��	<S�pe���`/.�`������<jIU���=l�97��ڼT���Q�	QC��a0��$G=��f���H֪K.,����,���iʊ�Wi�F�����$�ߊTw�tls�M�}K��y�p�޶��;�#I�{W�m]����՚؇�:Ô����(S�g>�	��{�fb�|�1���5M,Mܨ�g�C�'�=c�P>NE�pt����7G����|�e'>������,�n��}*1ֽ�I��_�C`��"��wDp��.��,�X5�GD,�����{�u��Ll�)��#X? ��V�	�r��.z�
����y&�ZJ>;������p,��է�;M*Q��W8�Elۡ8s�X˪��:jK�ZT��:d&r�p���첗��p���ѯ��6�J��l.��{�&O��ąI@���n�aSf��tD�����I�U5N�h?%vf��ZrD���S���g��o@�����C�]w������m|ڒ��q=?��^��E.��I�ؔ�Y�N��F}�g��)ԪK){nU� ����޵�5�W��V���+���E�ѿ6p��jK�(F\���!Fݯ�q�/��g����U9���L'�ο�i���ޓ�n����5PM<��c$�k��X��d�L�一���D8	�p����š2�"��S2W&G��|(T*)r�H��ǣ�����3�@�t} z�y��3�%�kz��:����5?����|��,3t�f����;��)8�R3���C�c��r� v��̴!F���V�U��dD>y�$UKM�������eG��B&�)�:gMzn�Q��H�6��"5�ld�<~d�S�Q��]��W�w�Q����]��d���Pw�c:���1���0P�4;G�0����l���C���ӓ�`��x�4��N�;Q�f�WI�8ˆ�S.�A��[�e�o2r"��R�]f/���5�����>���<�����˸�Sb��ٰ�-�P�Q��d�!I��dgݯ~��ϱ���u�m'8�-��b�����s��`�@�C�wc��H���D������x��M]�8�oҩ>B���J�����v�C&2�nS��X竩9���K�9-�h7��@�Y����GP�ƙ����a���rRT�����>`J��f��/��|�L�z>LP�F���� FR��2O؆�@L�6��P��j�����RX������XS�w�$p�`ks�r��*u�6��W=��NÚT��m�|2��͏���{��L=�~����,c�����52�����N�z/�a���r�	LR���M8ѥ�y�<YQ�Rql���~	�8񓧏�Zw��V������=l�!�9��%���T�gvZ���k���m\	���3b&!�8��#��'��b�͉dcA����>t4�l<���naB���ƵN�v�0� Rg�d$��Z�.j�5�M��Ӧ<��d�s�!1�翕� �_�u��(\���3��D���ҶLja�8WT����EZ�ϧ�a]b��O||�bt�n�[�&��/�}u���8�W�P4SQ��r�۬��N P����?@�w�Xg�?	�y_G��3�Ld9����g��nL�?;�q �.Vy����q��D3�U���҉T~yQ)@�ڳ#oЅ��5�F[��k�׆N�ej�ō��c�{xmZ�j��sM%8%��P������V�)x೤V}Ƹ�:��/m�7�ԊN�c�A�0�25�+��>#GoZ[��l��4�i�G��"�3BN�C!u�����j�&}ZIn_����A�O4T��[BiO�!V�Q�t��0������䇲��k����]'ܱ�)I��X�D��Ŷ���&���@�D�>��u蓅���a��ƌ��rlؕ�;axY� ��Kd`����d�)���{����ZM���0��Bnئٱ[�r�k.�.���W�;����hHB�L�.�p^p5�� h�|���X�?��1Y
 �t�������^e�P�w۞GBv�(ʬgD*�?u/�:$�Nb�7��g�o��R �$w�Uɤ3��qI!�E��I��YR´8Bbj��;��<7Y�h�B�ЄD��l?��ŕB�����
f�t43')�ޙ��̈́U`�C7T�p@u�j��L*j�(�I��!=�i%�:�]oB�N��0�T�z�O�!
�A��<��%d<Wo.cɕaY:P�4)o�|���տ��k��e�y՞s_yW�ix�w��b�#k��U�e�f�l����b��جX�:�;5�{�t<�~��[޿X�9,�fv]��A� ����V�!�vWV��Ȼ��B.И,#J-�Z��j={�l����`��aV xAȤ����i����Dikc������ry1j��8����_������Ja����7	R���7!����hVNQ�
�k*���b ����>�w �#XXdk�e�� =�<���K/���sح���^Z��>�:�E�l�LvG!#f�Gz/m��e���?H�����N
۸X��)*$�ha��&@4�b�^�}ny��G|M��c.L��e���qA��G���P�J��)&D�A�;Y{��g���y��W�d�: �2Yz}d|��Μ=ܙ��_R���)�QS\�W�����x����:V����Z��I���NPf��u�%9��{���(��b��oƉu�}m���z����O!����'���{bݿ�G9�ky.Y$�wJ����а���:�*��I"�21^�d	�W"U#S��͠N�;[i.�^����Bbq��S�c�³V�׋�D���
Qj�Ym�#>��l?�Ͽ�S�Z`:��;��/�Jf���L:��飈�t�nD���d�'a�^R���6bD�xJ����}�F�T�P��X���K�Qfu�-��4�����Т�i,ڪ��J��p��C�񖙎
�;*�US��Yr�N����(�cw���*�a��#��t]<�0٬�lD�Zo��5��?�A�;��P{ $Z��pq_Ӧy�d��NH����S#�	S����p�d����F���������a/ny<�E;��<�yn�z"&aD���/6d��E���9�T���U��'�.��e�2+�Y��٤I��]�:6�[V���֤�3j�,0�f��`;1޲p��V��B��4��D����o�݋��S�E���G� �%��Y:ZZ�����5MF;|?i�����Y��Ub�l��r�f�~^D��n�x/|��f�����Js�Da����h16�9��{���cΗ^�M���!l��Q����@�ẗ́�C��?7ήb��j���$�W9���%��.$ޛ�D�D+���󼩚�לc�����(W�q��vԞ��OLk�4�~�;�n�s�巊��;^,��y^��L��+B��S�+��j��H�+9�6s+ds�tJ�;��v/F˘�8��XW^���~���Q �)K�(��==��k��Bv�i��Nj�~7�՚���\��r����Z6^e�4>�@'�ygdÃ�I;U�ۅ�\R�qj�������a<ĴFo<�_ꖡc�
߉��LEpzE����!@�ٻ�.�~�e�K+#�hZ��`��fc^��4�\��*��q6At������B� l��(Kqb�g�Z]��K����1Y&�2�+�Ո�����Qi'4�c'���XT�_�aCV��'^uP�{J6�f+.�7���06���y���ԃ����W=>�꺘�0���E�+��w|ܳ�u���
	��:ERy9Z��E]�I�v�phe�Z�:6�� �А���V��Vs��D4�K�NyǇN�o�����:	��"��Ā���6=��>.��m��Q�9h��u(��Z�Ja0|����6N<���̞v���E\���*l�G��	���r�%gF/b�����]����a�ޢ 34@NR�t`x;}Β7bP"� lu���֤;M�z"@��ȏo�Ad�/�pu�FE�G��?�s�|��] v5-9��y��i��N���E�^���y�{;��M��"7pA/yMt�w�0eO�x���1R	�E���mw:��r����t�s$lL~��(��n���GN6`נ�?L�/>O�_l��G{�IN�!f�:� �mp���6C��:]M�$��;l�)`��Z�,�8D"+�NbJH��@oÀ/ˌ?�����ӑ%��Vr:�¤�^x���� C�>��8`��O2;d?|����� LsL��Yb�ko!��Q�#��	��6��m���Z$�I^PjB��*���Y*ɘ_�����bݧp�(�,��-O<[p���b8,@2�+^�D�,��:8m4��y��N����ѽ���ҹ�B�(����_���=��3�z� ����
Y�
����H��	@���jh}۶�rg5�O�2��1\�����b]���0m�7>�ŗ�e�o��+��
������?s5�Pq�X�fZ.�;zBb#��TI6Gz^�0P81�kbt ��z+�#�{Am#�&��QO����O�+�E� +{^�t�\$$���(2n"0JE�<���q��O%-�6NZ#���U����V&{χ�!d9�GPz�pKW(JQ�����ޔڡ��d/����p̅����%�oqT}��'�\�F����z���!.-+>�FL��I��"���g�~����Dxp�)���]�����O�v��AV�h"�3!IByT�Ql�|���i+�p܉���w������f���ߜE��?��f1䠨��)�����l�0اWL0շ��s-PF��Mx�C�w|�1�*��x�i-1m���F��g��M��x��15� �x��уZ�t�h�5���w���Fp!uAqQ�8B+J�Jq����0�G��,�/[���~BA��s��]������dr��#^7{�OՅ�2��1UF�9�W��7Un�W�3���#°2�)^��Z�o�Fǫ۠;�lX2'���F�L~,�@���U�i���Th�K��9C�M3�\�=}s���T0����fO���,�un�V!kP��H���U�b�Yԣ��Ȃp����'!86z�G~�>T�i�l��Z���E�*�e��u>�#R�B���~�B���']��%���t�rlcO�w���fp��V�@a��Q7CӪ���<������*�P��ۺuj�*]�P���7��.L+��)s��?��J�A9��'��QǍ	�z�c�C�cY'���m��v�[Zd��.�s(��"�l�&Y��n9�0'���f�)��0a���%��V&�Wwb���^7�q�����;h���v�3��9��u�}}��+�GD =�I���9#� O�W�nIAЍ�9��cx?R�
d���Z\!
�G�8���YKo�AV�2�ƿ� a���¼@ϡ��:�C��E@`2֗�3�.5������b�7X>��M�/�284��Kx"M�z����1Vi�w�������ZM�X Q�a�L�$:Y���y�vX��ae��K�n�d��æqňZ�:/Q���E�G�2��o��e�Q�p�;W�z���[rAHp�H	��DO8yX��0Ț���i>V�������x�fS&"�)��D3����GMy�cL0;p�3n�A"K�l�������I�D�/��=�᫙�*���]J9��c*�t`����6{bs�L@+�zH9R"8E����#�<�0�\ﾳEr<E������!��Yʪi�����Z���04�Τ�U:w}Ae�đT���*��/��g�}�����i)���� 'k��>߀�ٰ�q��ƵƄ_�����`u�B�g�k���z��qG����يح�|�����*�N����n�G��׉6�5כZ�>ߩ
_9��>�v��XgC1[a;���;7�E4���<H����N�@���D�]�3�i�$�U볂-�� W�΅����lH��L��$t��V?�CT��Gsѯ���!XHx��X�X�>������x���9	'�@:�@�qk���׀����	�_�U�	)�۲_�9�+��7�}�=�m.zSDћ`�R"2���������v��@*�%����`^^S���{��	ኬuM��(�8pǄ/!"j�,�`�Zmx^#{�Ɔ�Qs�����u[I�<o$|�{�ZMɞ5w�1:��ri|��7�=ޱP1�6qn$]t�R��`�B���3��K�|�Vn�)DE��н���]�B�ڦ�Ax,+�aO)h�UHC���(��L� ��$gM �AA��?C׌
� w��(M�[�2nA�����0�=
�Q�9��})T5�4 �����;F�V�SK*��R�?Kh���GٰW{B��O���7���Ǉ,��ї�I��9[
97/(�+�yF�p�W����g���vj��6&�\8Ъ܉��A�����@M���:�GpNd��m�cɻ*�N��o���bmMb���d;�MI�����,�I��C��k�x0�i��c�KzSH�?��
t?�P�厐ס�G�!���x���H�e+X���T�H�?�Ҫ��Y�d曁q�_�tɫb�y���~p:aSO<��o�[��'�P�#�[d�"�'��p�����	>�L��-�+,����:v����!�p�d2�5-Tcw@�f�Tu�yN���/����6�D0������w����@uS"�/j�7�M%���MO�T�͹��&��,�f��>"��ʥ[�w� (و��+Y��v
A��J��q�^����%�ܡ�� `ܗ�i!4,���U����
�K+"�B��3��h)��Y�UDڭ�m��5Y��Q�t2$ɩ��S�2Ƹ��;�ק`*�
NJ�c{cDYm��#����i�mH�t�`��?%�D龀���*��r-��ͯ��j�����g��~V�62�f�9v�20����[��?-$�ͤ��(*����w�2�q��ϼr��rup``��
���y����r�̜�xA�g'��C?l��LH.��P�DG�ΐ}�L���ӍLa}'Tp��N)C��yۃ�s��aE�_$%J]���3��p���aMՅ��^ n����W�X��XH�]��
n/B ְ�X`�	�u�� ģ��oե� $�'�
X̃w��[߆�c��E����k`�Q��Ӱ�?b��|���6��!��\i_$�;Eu�>R{�i"l�5���t�`��Ӭ����F�޵R�pP�D�9�Z��!�0�Cp��rӨ|I�
]�5%�M
n{S��m������|> �>�/����K5FߨZx����7�H�;����q�|�s�3���E���'�<�1<�
���dIg��$֢|i>K^<���^��<|2��Yb[�~��j36{$[:�d�$ho�]�J��2�Jš�a6���t���wa���) k�W���/���s�\�JEt����8�S��Y��{��]�:pf�$����`��3����R>���]_3d����"���'����%� F���=Vd�$]� ��JEF�?}U�]�7Ό0�`��\�P�ǔ6�������28�n��w�R���	�N���jD�����?�,5�ٕ)J�:y�h�������EEZN)Iv�6*����+ݮ�X���`��$#9QG�������C7�?��9�WO[oC�u젒�}E����8�7���%dX�a�ԗW�����H?�*�5ӂA������4Z������j��Ϋ�2/. �f�g1}x
)�I��\޹ݜ�y�6��F�lBI�����E���v��X�u[Ƽ�gx�˓��V�; d�	��#M(���9����B�!���<F|����P�F`F�����֬�FLSo�9���7�ؑ۹Ա�a�S#vt���'I#SD���	PG�K?+��ۖE��*M5� ��sb�'�P&�}{N�g�-S���)#�9��������7�p�OQ?nR�OUclH���d�+ڱ����
�"�,2^�8s?u���Z�j_�`�k�e��=%�}r�Zl�/���HXR��]��;	<���eL�qd���'����j�n�2F�uJ�hM<{�b�,|Ԍ0m3�r�:�m�P��z�`��±�^�%�ko��\���5K@��xD�L��d_*Pc�1t�7��}��w)�����#��JIE�s.5�M���y�N55���|D���_"��7��;ǽ��b�}>���;M#ibZ�>�ay�G	�ˡ7r���� {��������z�Ma��F2`~@�l�m�'�S9��T�.΃S�ڥx�,ꅫ,�k��*m0�����|@N�.��+��I��(��d��d��7Nk�vf~u��e[V7���t�k���BSwl�
�I�iZ/[�x��֎!4 \ps��D	�4�Nh�y'���|µن���B́�T��9�*˶@};����s�̠g'!J$���p�>:��Cv�c�����ex��6+'��I-�b^�D�^�y���n6�2�5oA��ǿ671*c��!n�M�g,O��� :@�����[	��6W��7��OQWq�(�.��t$���R�<qͤ��}��۴j�i�K
py�[\��E�v2g�=�&�0�'����%�n@g�����Q�Nn��AE?\^ĳ�`��� L��M�_��[���Ϫ�:wO-}�Ɣ��:��>7y�Bز���]l�HV~�����YnǮ�Stf|��(~!RGLa~H�IҤ�D�k �#}V���
9+$1�Nx3d;Bd-Wv�NƄ9&����RD D	 E��Q�5 ӌ�l�����6�U�ʟ�۝���5+Pv�$N���	�%���us�3u�Q�ߑm��_��5�'w�x��a~\��W��]�&�4�ر�Ӄr��.���"0���l$�`5��������_��=9�
�U!Yr)�Vu�Ɯ�!���"���z��a�'���l�ռ�ZN�͑m�-�.z����u��A)Q��؅u�|��������$J	K$\. ��
��S//��[<�_fV�Z����%��w���
I���,=a�@%�\��?��p��u�/D����r�s^ؽ��ε7�v���Q5B��5�VB0]�w�a�����EM�L(?� ���p�?Q�Ak��5�ֲ�:
��a�c=��+������r^S ��)������k�~�KޘEJ*��0����f�l��>U;l�#�fX��t�^s�n�H��}ٓ�nvHn����~lV���V��tNI�?E�T8��`�賡�uNE$�WӔ��\�$(5ؓriW��IV( J��O.?�3y��&�t��[Y� ��U��8K��<��KE"��a���,8'��j'݈a�ǔ�m���h�[2�[�����s�H�kj����o���`8ĥBJ�)|*G 1�q ���1�	��&D�j��؄b�ϛ;�Faχ�o#i���L���ҋ�XO�%�j��4�?,c�=�y+�ϻ�l��w���6T�D<	�����'�VD�g�I�z�U�\X��<.^=3[JI�5TTֽwZ�&R!�SF����Q�hb9��f]�8�]ꎔ�Aѕ�q(1p{�m�c��ؠ~J��_���(��� Rɚ	�b��߼����\�|���Wଃ����$��ǧ��*2�e��M�y�`FBA��r�LD�
�U}`98l������އpZ�X����Ә����nۄQI�\#���b���|��2.PZ���
���k%n�_�%~�/�dw�Ĳ$�`P�� ��?�'#�T�&(S�8+|V7����VIh���2����� al�(�5�}�
��+��o�u��/���}(�e_b��\K�3Obw) .�A穢�#�l��Ϙ1�k�
ĵ����������+qp�FM>-�^�n&��� ZDH
-��7�~5fr��f���-�l���Ӛ?����bT���F��}bm�l6���W���0UI�E���4Р��ղP�Buq��=c�s���#��xx�(��PV�,᙮Sk���;���x�?���^>.�U���y���=O��+QcA��:���� ����f��:'��k�g�����d�f��!�;���ձ>�)��r{��n�T'H��0�)o�4g��m�/�A���x�W�6��<�'Ů%V�C�$�'Sf%.��tk�K��T����cI�䳊���j8�i��LWµ�&���uP�nF�e����5N�,�:�Q3��r����X�����U�'�Xu&��&��<������:3ו��d�O����s��ؙK:�C�c8=`IS�i�^�Y��u�v���#���ʞnv�( o�J�yTB^��OUz�#˙1����m9����*�K ]Dv����t�cU�:��"t�D4�������mڕ�'���Ny�`,?�Rj�K�*3	:�fYY�)�gڅPOt�R���#�Ƣ
�I�mA�<�RDxe�iI�.��=q�ѝ4��_
��@-�'�,n���E4��o@G�'����auM{���U�`L��v��
s]炴�Il�A�ȂXK��dKk�W�oE�ФI=Eݑ$'k�������\BpBi�X�8T�}��o�c댏 <���U�[�lr�"�͑A�?QJJ�b��m3W2I�Z$���1�n��c���a���>�>2˪�u�M�$�6_�qV���v�O ]|V�K�_g��1��
�lI�=h�2��_����̄S�_��&�ZE���1l�_	n^F�x �d�ԉ��#��.1H3��o�J6?�������w0��#�>Ol��a�3��rM�sY6v(��Ry��QQ�вB��T�����e:���	Jf�	ݰӖ�Z�,�b��э=z��ifZ`hU1c��Ԅ�4��A��%&�/�apѿ���4D! ȷ��\QU�Y��*�V�8jG" �
����E������g�o���^�t�:t�|7V;���*�۪n4���LN��F���}	Qb�(��??���M�i�)���VQ?-'����h���խ��4��.7Nˇ���Ch�UhGNfx��^2�����H�A���J�q��8'E�،�$0_�em���\u�����&_7�w��`����Ϡ���_PPr9*R�K6'����K�d���w.Aݹ.bXSƅ�� ��YNDb�]����qP�t:��-��h��h:)#fiK�3���;bs5��M[�r���g*����	p�ߦ:q�ʾw���P������XkQl�{*/
Y(H]˯�du�\�����N�h�[�]�3~���?�-�sJ��/����j����3�s�}f�*ܳ��^��,![��.�cX�P�oC����o��Z�f�egC�MW�K \i:k,�Tg���$Pȳ�ѿ���$�ǻum.�F���&G�R�Ge*������8���Ἠ�i�3@���F2*�A�����u�����,��C����w��(��|C�@\R�[C�8�V���1���]�<�Й;�
9Ƹ��T�k��jP��K�έ"�1�$4��ToIeD��qT>�KZ��h�T���G�ziꁙ��D��4�{ ��q�Y���gl4SHXW�^�� {�Nz��b�붯�+���^+X�R��8אM����*c����h�6v;S4���^��QQ���7�h�1����;K�R���V�뱊�a�:���(㽭�����{8t���d�$�S���6K\ABE�y� ��w?������T�lI��D+`�Q�q�`�웣��q���LKR_%(Tc�Y�0�_���= b���.��}`��
7�6$0ui�餉���\�k�XhHl-��ynq���i)�J�C����7܀���[ub|W�����Ϩ8������&��'������9X� ��	o��F����&#���y�/�^��=�Ǳ��m#{��gͩ�ڷ;��M���Te`m�n)۔&>F;9��)S���4�IΉ��M�]qrry�l�F����}�%�2�Hz��IYPb�B?�s��Hs���]\>?aKE�a�.�>Y�,���,�n�P�8=�b6n1�؀R���zgI�uI� .��H�۪Y��*�����@�쟓o�K�Ol��c7Ɋ
%�#O��[���p�{�Y\�%�3������:w�j�d���<v����O.��`iEW	%���y�ܱ���:4���Aޞ+��Vt���|�ƭe�w0uӱ~�m"�J}�`��,�'>.i=��"x0�2�$�����iU^3��l ��!Z�#&���$#�Z�o�QIn������~*�t�m�jd/��J�G9��B�Nf4K0�{P4s�%,[E\<PPĊk��ۈ!�bF5�z���{�(���O 9|�����?ܞ7Rw��������d�����`�cu��fe���%��z+��
<S,rM��=X7*?��6�f�?[�M��#f�Y�T�E��6�q}%���֦�h,}�&�����S|��"���X���g�It��_��4G��3��#jq��z�U]���r]/���4�V6����(*�< �����Ud-T�G��� �IlU
���P-H5�1}����e74nl��ਜ਼��iU������|��F _K03�'����� L�k~�Z�N��a�Ѝ��ᚩ�G����P?3*�h��d��g�碭���C���xHp�h�~�� ��3��<,S�p�~��;�t�μ+
X)�gR,+�o�j�2��7 �;hyÅ5��\}ޤE���]|&��ULp���������~�P��g�z����J6m�T.vB�J+ڝZ�p��XW$���~�X�0?PYGF��A�@��l��3`����{����>ٞ1)̖M.�>MinQ
m��T�臇���������M�,e��l�^m���H@�)��%�g9�Aq�:g��J ��`E�A3�E߂��E�. ��>$]Ń�ǿ���>/�Ki��?�*ˊ��!A�c�f"X�Zʬ�Q����@ej���sꐐ)�o��w�4�O���Lz�/�L'�k��X��<��t�Ȭ����RhɃ>�����Z�N��Ϳ��}��$�q|b�yw����r�� � �%�!}�%3W��A�[��j�����'Z2��	�N���p�M�ۊ=�2;.��S�����[=����S�¯�n˶}
tFQ tg�E',ͣb
ʺ�=�}���s.�4 {�o����k�bЮ�\� �N?���jE$Kw�Cڟ�`����y�b����)\�x���T��*���]���#��;"җ��ȣ���:�fj��5s��S�_�=�`� ���J>,��D���c��$��fa��^��Tu�c�u����N"���T����Qé%Hgm��������R\�X����H��kc'{�t(J]���:�cE7�r�1'��ⴔ}�E|��cU걃�k����1L����n�����\;�e�	ؐ�+e�_Ԝ����
��Ϥ9�-���U���ʂ��U��)׫f3.{���	/1�/���p�����l�l�^'3����{b�|@DA%oB��(���b=!���lm\Y����<�W���I����<`o!W)\<+e^{U��,V�`�֙�v!��c��j�ZC�㞅�^F-�o����zh��A��iw<G����P�#UV1-yM�"� ar�W�o(e�����֊������>=g�>�ya���H6pЎ�/]�~�k :�`йn�H!;�d�iX��]q#1۠k2ͧ[���w����?�a)�wo��[l%����aV�i�s4�;�����]�J�pK�Ν�_w����m�5?��r�-��ƴ9?�n?�&���v��<�� ^��M����J.<ZӋ�̅���䰙;fw8�Q�	� ��ru�Hz�P�yFrd�W��M��Ͽ�*�:�N��a6�SeM�u]4-8���G�' �������q|!;ꣴR��]c�����_�)�u�e�]�+p'�n��v�$�ˠ�[�?��J&,(�9�����Vv� �y����g0|�%�d����{B���@�qn�4���@��y�?G^�����B�ܟ��#�7P�1�U��/8�ѹ�TMü�Y��;
\��������]�(j�5��_a!���$��s����Sh��m$p�h���U����|�,'M�};�t<e��x,Ó+���PM=�Lyٺ.��n���8�O������_����oM��Vҡ����RI�ǡ�8�]&� R�5}���g��?)�T�v(?�Q��������a��0���ao���.$O��j���@3XqYy){ː�
��V��1��g���fk�^+����D1�Y�0~���b��G�,�F�E�x����&�L�C��K����T9�ʺ�.�k���CM��"��?�8�E"ٷ	�ɢ����]H85�`ת(�1&LJ�>��.�������N{�W4y�q��1
����в<J��F��?T�l-�h HY:?��Z+Oǃ%$���<�Q��5!˜�L��f��[ S5H�%^I�n�l
����[��^�Z
��?�2���hc;4�k�RI	@O��j���.3�?���a?3H^�����I4M����e�Rpo[	�@�Wb����B��:�HDW"Ř%}L�x�[�mY�,KH�HT�{ohD<����ؓ��8�ό�Fs��N���/�)/l/��6{�?_�u���bJ����_�����4��)W5��֗m>�#L�/ʥۅb�P���L�*��E�/�V��Y�K��Q�A���.�~T��&H-�?t9�y��g}������C��u����%�+"D1?��yz_;Ҕ9��u��zb�;t`�yJ'�*�MM�;sӣ����:�a%-��@Im��S�dO�/	�6�Nw�cA�&����2P�ol����o��Ç�A<�k��t��"33�K`�G� ؓ�Ј?�Ƕ��E
 YTj�PSwx��;�	�����F^?�w
���g��<x<]�Jt�ΦH�ԞU�#�o��eަ���ȯ��Rj�(��Ap��(J*��.O�Z�z^}Y�jb��aWi+�Y��+�oq�_z�Պ�dԪ�i�l���V�r��{z�{���)�-/�ؙ�0's¥���y���p�^�ؘ6��T����GTP���[r*+�^�p�2�DvtfÄ���:��:���{�h��jfGc�"���Ys׼Jh�����t̪.�qy���60ZÐ�9pe�n�|��1//������A牾ӟ� �1����K�:��lC��C�*-�x��i�NNد�D�0��hK��� �p��L9����&9�R�մ��J����yF0�?��:��6��d������B��#��E��MJ��v���ݟ�'�Hg�'x��a���\�#]��V��\��H1��`�1�:�81�e�H��$�ZKJ��� g��v�M��3���J)���sfp�c�:V���sO9���"�(��'�����X9��$���G��1�����+�N��u���iBʯ���7�B.MP�٥��5ة�E��~�C���L��f���o��y���|� ,�%�����ɠ*�7Q$��DkI5;|ha��-<Wj=��S?�������w�\���bqn���4�4�\��
���e�j��\��Z;Q�i�u����<aEt���-	FHO@~^�?%�����j�A�N�b4��Μy^���wQ�3�I[L}ˠ;�Ow�j�駆P��V��Cf��Zsў:��j舊�2���XeW:`8�g�F��R7w^=��I�@�����L٠�m��M-����)��T-�ٴv���JV�.�$�Il��L�F�2�#@K�z����`9�S��b�x2wũ�g�v�I�I���\95��b�h�1�we�9�]@�^�տ)}��>��[7�d�u�ߣ�������̞�'���ES��A�V(p���=SQ�F0�U)�[%����$�!�۹X�q8?"g^�6����g ��̓�9 R�9�.�@+��R�z ɔ�F�m��;� �zx�u���X��ZF��Z)��	�ۣHځĪ�12uOE<��O�9I���/	�
s�U�����}�c�
#��λ��P�龚m��&��7���Ug,�d���U�eO�T�4ٯS�0P՝k������A��*%�ѕ�F�4*�z��A1+�'%���Xa��hnu!�>�X�(�6��p���O�u�r��yz��E<f�L�1����|�����y[�Χ��9�Ht&�a�$��tC�K�;�YMFi�-�\%�*�a�(d｝�Z�zD���
%�⪕��m&���4V�.�Q������.�<��ҚC f��PM�]7�$~�iԳ�]��]'{�D�1��}a�����򠲝B��]�W���_3�	�JVC�O���b��	�9�n�Q��l�n[�o?��܉o������a�fY�t�bJ��K8��_��v�O:�Ƒ��iJ����|J �L�r�ߞ�Q� ��
��L�&�.�6����𯋀׫��?%^/����]�>_ņ��!O���l�U�/dT n�4����/-K����|�i�	����يh��VP$���|��~�e/n܉D�RGa#��,?�b����v�:��#�->R��؃�G	�{uh^���60Ӻ��W���Y�Qd}�2���JCZ��S��1�F� ��6��$��K�kp./�y�7ڔM�Q�d ,��[��* ��Q��j���� Tu=҆f��;��j�j�A��'�>�Xi�3��ːM[��ڪ����+���P@�0m*Iw<�}���D�7�����sVR8��2�{��r�f�%�v��F0���_e��V�P.�EB�^,i!̈0Fu�Q(���d�`f.��L���[��,wW}�!���r[�S{��Qڸ���:JH�������@[���bSR��p
޳ҫP�,
S`Q��ʞ�`���e������+�d�i>���-��V���9��xc
��i�c�LJ��B���gґ8�N���D��QɆ�{����1��}��]���������}ˆ��`�
 ��Arg��w(�d��Y�[7���;���-ᘿ�[���O�do��6�� �k8�%ys��>\ч[8�ce�N�!�2F�~mt�ʍj�geq�̓�nr���;��t�����Xm��M�t}�<��S �+�����ȧ��Z`�P7~��T� ]�	gb[8V�~����*���=�N�E��҄ZR�D@�s7co���r;S�DC΄Q��8�C�}��3��	������?��88�`�h��~�5�z�WT�弋fi|�ۺ'������+CL4?���'��׾��W!�ˑing��gS��	Șy��n+�y�^Ut��W^�~!C��'�d�����`���-��:.K�l�X�N�!�����j;CO�{G���V@�7���gM�"���츭Bȳv�BLeDhJc*x^]&�i7��9Z��/+d)�������0p�c�PT)���U��r{r�n�H��
�b��Aŷ'�誷����=��섰u�n�i��[@�1�Y��Ln�>Wm�jT� gL>�T��~�4�{�j�����0�O��o��������خR)���ݬ�L���rI�r�̚35��"���ʦ� ����0b��Yxs�����'�Ď���Je�+Y�T�����Y�	U����k��F�4��������݊N1��߇���;����"sΜ��Tl0��-|��>Zv�y��E��\����[}�����- �\Ւ��d��/�e��n�k��$����(��Ʋ� �V�� �"�H_��y>F�j/3��l	k0̲Xi ��y,��佘� 浵 ��%4�M�������İ�t�j�N����a��IN��%d�B\F�%e$iQ!�����Mվ����W�n��� R�[*�Vy֕�/쫕���?��E�EhϾf����}�^�L��ɄB�(�3Ʉ����?^�!�c<���]��C�����]s/�7����Q�E���)�@������QSP1�	�𯌠�����ds���d�dI��t�JCzd_���u�%���@~6����m��������S�b�J�wSc�QF�����"1Pe��h���i�Ȅp���=Z��3�{R7t�.�S4o�Q�I�G��oX�v�G�R~���(v-��4���[�uI�0#�-����j�	�|X�� �R�f�Y� :Gzڻ1�l�u�W��+��Ŵ��.ZO�o�7���Ĳc(�J�^3�L���%�j��==K�h�������t��}ơ������h�����CN�,c�F��>2Si���V������
���1��\�v�(,25T��_��/;n���k!>��M���b�F}��xzW�����&�dV�u��{S�&΁�r~���,�>�VT-�Ue���NR3;�ov&����Q5�l�z��ͪq�!hb� U�O(dS|��4��v�6����.G�*"c�����b)��*�k�K#���l��Hn�9�DM��{����[u�{mx����p#9 epad;�崲�a��.cx�&=O!_}�$�ۖ�E�Z�!�13@����`b����P_R�ec��NJ����)��5�R��Ԥ-������喭�r��~%�AW�Qd��l�Ki�1��.)��s���}��������J4�̏i��(.�ߒ?L�+t����v�|��g���-9�� �4HAb�M��V{Gl�+!N�(�ӤR�Q<�F:�����ob�r����/�v��rs72lw�4�W��yr��g̈́~cjʾ�-�(�e��g_ �E%;�LS)���gF{o��i���W�6z"^׆������{�KC�<����9������B>Y���J��?�e�z��H�9:���=�l��:��MQW���5�B�z�Tm|���d��QZ#�O��/L{P���g%a�F�}8���PohMkc�2�^�h�T���E���an�X􌈨�Jv���F��(426xfٰ���5]zJP�t����t�������ׄ��O#tT����aBq��w*�%TS�9��@��K�dѪ���A����\�bX�.�V��G����uu�:ՀHC�1�~MH>�*�����,��8��(3Iη2��ւm�sC1}o��H�mD�5�<ܩJ�?�Fe�!�M�q�ŹiD�;�
�	�.��/��*��d�G�qe�>e�r�� �/_f��ZA�^�fn|��,�e�:�8�Ahk�eg�A�e��Xe�.�A}��'OmYS��$��>��ٰ�|�o�d��Q��>�Bv�u��o�׺T?w%՘Ԅ@c!�Q<V+�6	��8|���%/$�r��&�
�\�-Mҁ��ޭw��﷔����g���i�^�
i�G��l��{���6Kף�� �q|SP�tP!���%�;��bd�9-����ԟ�&��y�jq)���S8jn�	^��/`�q����
Y;45Ћ?r�zËqh~��D &/�h�qn~���g�!Aĳ9� D�XS�7/,�����P=�k�Hz����ut��[��{>J�v\71�u2A��'�b{�X�{:	��N:t�Mud�
��6�-�+�]e�� s�n�O��g��A�ggZ] m��J��!�~�*�j��g:���f�.����9�����1J��[X:�9�`s�o-��t�
�As�_�I\��?�i	�8�R܆����Fj
��r���n��P�K�,w�%B���#�9��j��MkQG��(�6���0	��U��������~Ϝ��f#���(���$�Ǝ�������ZI8? yO�2�0-ޖ��`o����	J^*#")g��ǣp�z�@��0�X�#V�G�yW/�h���sD����c$��VBi
�SF[�p5��d�ޏh��y7��W�$�(�j����꿯��0�/��#��Y�i$��>��*Y�<g풣�u��6��S�6�Hӵ�F�u�z9t|�F�
,�q%C�UU�$��Z�s$XR�HC|�����V�Ӟ�)F����<��Y��t��]华��8�Y[�bOs ��=���d�"+K�(?�p�gZ�u��� ϑ��+ϪK2_+w0�T�3�$LӮa���K'5R�ⓚhSJ���a����/�����X�C�H5�	�M�(��A*Mb.�˦u;;+�⢨�)�G.���#��?�>�DN'�>�ǋ.)~��)Qy%���^ZN��$;.Z��%�?Li-������!w�� V+S~E�s�����'yv�F�w��ׅ4�x�T�zuK�+���4�[<ƍ�����V-��^�R��=��*v;#�?��-$#��[�bvyl�0	�!Y0�0´��2���ǽ^5�5Uy���T����!��C��1P��(9��Rdk�9ҩkm��ҁO1t�R��_�M�jB%�����( �*�揕l��h�=�Sx����6�2�E7Q�g�<qd��g[ki�µ�h��cvw�P�I��-(�R8Q���rͪ�V��d5�p����;"�9��	W����	�:����|��Ӽ�~�x�0���@�eڪ���1�5h����aQa���5�x�NF�`�ӽ��R�����B�Iӻ���Wo�Q�Jn���^���͓5$P��Se��h�H�[/Ͻjj����N��I�-�`��� ��6H�JL��p��0MN4�:����	��%k;y�`�^��r��/�)jx��g�7���0�m�$^2�� >oo���y��,�ǯ�����(K	�>Nrf�q���V����1۵Qq݃-y�vQ�ґ�+�f�E�ց������U��(�6�����Lyz"�,�r���<�T9�K���gÎF,%�&�f�W���;��a�>z
���Z�&��hz&�Xպ�Aj^W�&7�t�V�K��/u�j�mK;�#<ké|�->��Fc�����z��Ӗ����������[�?�k����(��{�8T���Zc�ֈr��H�JJ+Z��Y��a$�w���Z��u݈u�R]�؈q���޺GH@�"�LY<Ԓ��E�}f���'b:du2bt�&�6nb�Z%�'V�擂MFjM�#�ϴ��;��n=ܓGQ�p��3�cr�I���+u""����ujXr�����)ǚ+g���?4�U����/A�1�@�OC�"S?��L6��R�����_�B��>���O�V�s1��V%�l��%>7��C����6<o{�'���39k��ߧ���H yU�VƎ�E/��*��d4&��/i4�K���Qѿ1���ک\_�������R�)M�OfI"���I})���&*���f��5��e=t��##ğ�{K��Ԧ�_�\ѓ��Te��w�1�jd�rne�W�$���`�Py��Ḡ)�y�]2-��Hf�Q����B��g�Ɲ�v���q�ǀ"!!K�5�C��#%b���*�y~�rm�<A�%�~�_Cc�8���n�=&��n/��2H�B格"�#�4�o&���%�̀ɤ��x�%>	��ɹ��E�l�(9�V��s!��#���֔�|�X]��,}-�v�,�X��I�G \���=���}�WJ��ˢT!u�F&�V�u���d�d�*�7M,��
��#�M��D��A���#=�ʷ4d��Z��SK�r4���´z�t<�]@��Twnd���AE�Q���1���G�9�`�$%��|ӟ~��v�(�����h�4yiwu�"��,|�GŔ�-�A+��;&��FՓsQN9���z̎��4&�YTJ�\��֔���rL�'W:�&�?���v��:7�m���D7��.���xZe]����iu��O������ּ-�UqH�\���Pn��B���`���($������^��'�&��0�?L?����w�(J����lj-��0X��+ò�W?��9�΃
}L("���z¿t\Y.��0�p���3��!��b�bz9�/�W��.@����G�0c����S<��Ž���勒��,��P�2v���Y�IܧƆ$D��3�_�����z/r_�$�Xhe[e&��X�P7C�w���jF��H>g�~�;k��-YՍQc��2�|:����n̚P��?�7�s����O�l6-��/�6���CZ��A$c8�ݑ�	Z��
j��!����ۍXV�?�� � 	��JI���,��!l�X.DĩR�U'������|�C���2hD��6���B,K��	q���D���F�>Ib��7z�7d��8���)AW�PiD��3tjx�R{�r�E	�����n�3�p��JE���D�q]p�IڕMb>t��MH�?L4`������|ėq��3�[i�²���B��(��;%��,�)��h4�^��}qx��!��^��y揽���7�<�ȯ9�W�I`�Gp��Y�>��R�Q�|~J@"%>5xB�%���� "���,�����E��k�֞�b���c(Ri���%(E�lа�\���m�q .�3�QE�Yq�"veI���D!�I�~md��@��=�A��,���q2�J�|����ns��|U��푛?@E����s��_�J�[1��k6Lz�Zdr,�'W�5��I��UV�A�u�_��r�|^�<2Y��I�`ʹ��v������łp��0�,\�%�N��K��5ػ�7��%�~[Daih��f
�nd�6�r���F�#�0~�&�B^��og��Uf�Z~mPi�?�[��$C����=4{�����BT�BnSK����ִtp��F��)X��tԢr�5��]�ժB(ԇJ�ah#��-&�7H\�������m	�,8Q���*�%Է���x,�"��<̂^��N�P�1*������%l�y�/g���&ZP �ѵf���`[K������>�߃�ٚH�%<qU���ϝ�K$J. P��<5~������u�V�L)�h�%J�g4��+�	A7�|�W3Q�A[-�e�f*ذ�o��E�+/E�w��ulX磚aZ��-���@����9��-�={��p����3W�*%��❮��?a�Ȃ2�-��:L��H�iN��`�le>mE�#��hR����]���t�/����?���8�)���9P	Y'����	Y,	�$(���[5�]��� eKT2�B^2AA.��~V�窧���s�Fӈ�-���/��B_������s�����ss�$��T,���8��
�h	�o{�uKX1�2;$wO]�he��ې�b�j�zÿ�]!�7�S�N���,WP/�M���=��Pk�>�Hz����(J��8�njC[(�4w�*�um��>������T$'��%"�~��1 �w�����h[��aS��Xq��"k/h��(xd�(˒�.�Ŝ��T�1�R�i��Zi�����wFg�Q�#wPr��Vc'��{���O'$��8ݪ2�V���tS�G!����A��f��IH��5�O����xP,`|p���~;���G�?m1l�@s�j�Q�\������x�X�%c�lֆ~]\)����_��n� �
���Ȓ�7\���!�l�MԱ��t��a�NM!���-q"��N	
@���$5�����g�������[�#�_H�]�rf��!�Jo
�2����9�B�r�G�h�zE�]�����]°,^��ӱ1[�8T���ks�2c����u�r���{�� o��Qb{�a�޽���R���屍[���=6}Է3\nL�o"Z -�O(��6�|�w���4wm.�<�$�l�P�<.,Yn���V�U�E�s�� l�Z���zU+v(�fywbeC�?�N����oC6�A��fk�͈���}^�s)�n5���H1�XFK�{hE�wh�L3����0Lc\�-��+��ن�l�9�.�������Ί�o�1nǓmل�~�T��@g���pЃ�y��.��,qi����I�ѣu����uSG�R� ��VI�_��^�����I�:5�b�*ʧ�~��&"�^	W([�p�PH���fT��=��d�?[�N����;�nzrc�ZSY3�1�+r������jx�P8���5d=�6y�A�$�M��{��-̋�-.?��Y�7-y1�P,��}�Gf;Fd��nD�x�ປβ���X��~��r5U��Xj�]?�m޼�]�+�)��m$�=������h�=+[`c�3������n��+�9���K��J-�9�h�蝦V������'�sF'u���3W{���Ӎ�Fl
-ih��|���+�������00C�����U����i�+��>��݌|���7��!K�O?��;���e���Y�'���Q�'�c�ھD��N���K���U>+c�B��U�̲L�cc��^�5s#J�Pdc�-L<�3y�fa/��88��v5������~�b�n�wZ���ܑtb �V�f A�w����e����J)fp	ܪ_��4��Ӥ���\��Vb?@�GhW��+/7��l��#�1�c�u���s�4�&Y�i�E�55:�ɐ4&�<8ӻ�5�nt1���`Ή�e�Ir��b��2o�蝎�+��q&�_d��Sj�]�~��;_k��?W�&����J���;Eb��}��
�?�w�Kj+�Lz3m�w{����!�������&
�޸A�N<ҿX?�Q�Ie�.|��MOr��G����!u?��`R؏�ym�O�(6�uFJ~'�#H��6��l��ն"�mM�q�%��� �.7ԍ�:�a`� n�ȍ%���] �#t�%
���?HJM�A2m�r����hY�e��/�D�w=��]T��V�}��CgJ@���߿N;�V��rp�Os��'s5��ЙZ�M��ep�z}L?^�r3v��Ȧ6���]� ySú�@������Ux"��rڕ/&�(b�B�r�1._t~���T�PMq�^4�����t� ;�3FE�i�h.������"�0�9�.���n�<���︭�P6��rvR)a�ȼM�w���ր�+�!�K�?�ׄ���ڨ;eJ�솟����T�6��$̷?__
x��(k���)�C�6����e����0�#G 1�w��f��)������V,2���\�4��7S�ِc���G�t\$SJ���e��08�ò�;4o�<�9l%�R�c��1@kٹ�N��^G�X~їݜ�%�>��FQv	b���g���Z��n\��t�*EmS+!����1RD�5\.�(�͢�oBYǸ��U �WV��H���srƢ,,�l� z���;�s���}2�z�[����C��K��j��	5�X�aI^����{#@������r�3��x����D��x��jy.�9�Z���V�׬[XV��e�eLwɈ�yկg�F�Q��tj
���u�~� ƀ�Pt�y61L��Q����&m�9c8��+�xլx02�����\��/���R&ZR�f�}θՒ�}@�u%+���"&E�s�fl����x�.\f�P���U��c�?�\oa;ާe%��,�`%�A����5p��S�麗w{IF_R?|�(M�ߨp�&��P�j�}�3.�t�?�P�:q&=�PO�I�Xԅ��oO���)u8|���u��qt�mיU�ԩ��ƥTt6�8�]�˾C*�DP���l�}� �E��.K�po?ň����BD>)��|���q;�ݘZ��%F�:d���p��i�Z�%["
���B����n>�v�ͯ�&�i_��a��h�x�������=�*�I��{?�#��x�#52G$���
L�8+�#+>[q���
2:��J��N�sϢ�6e��������1Hu�vf}�Ll{�4�xz����ޝxK"U�~�xO�)ܬ�?gdj7Ĳ��k��Bq}
%��9�1y��]�>��֍
�V%��m�nݨ@�ԙ4��_�)���YFAH�� T|,*�Z.�$ǀ�O7Yμ��n(��}�¡�ls�LiT���'�+n"݌���N��X��,ڷ!�_;>��܏AYs�k�}h�N�%5A�_mtk�
�u�Q�j\�B`(��<h�P]G��|~x�=~ե�������7��2˴�Z�/,�� Pb@޵�Z05�Xe����	��a���tn"_��	�U��5��[��x���lm+6�Yϕ�94-��=5ޒ\t3�{L���?�����Y]$��h��h�M�0�8�u������毎�2�hY.��z#'��t�k�YQ�\i�
���_"��O�&��4��+x����jP�s�k�֢�f�:sA�+2�<`�Jԕ;��ojPp�(S<r�E��%l��M[S��tRu���'���f���(s�sw��Q�97�H����_�������ɎU5r��yY�o"\�]��\�2�Tk�¢
�y�weI�a��Qmf�/-���5:ο!�>	6\��R����+d����Ƒ�W�}�y��CCڊ��WQ��t%Ȯͼ�ii��mָ<�IM�{�Y}�~��/R�d�o=C����ب7@��.���:���޾w��=�SuYZ:ʑ�(�y�׋d�הC�޾F�l?����` ޤ!{�2�+��n|?�0G��� 2Wأj ���j��"�J[���H�`ꉂߑU�EL6��G%=����ȨoD����O�g:Nx]�G�z ���c��U2/~�z��,��5ɫ]wk�f	�#�.s����n�Z"�t+�i}.)����h�!�|^�h¢��_��Ra�u8��=n}n��BTM�@��]Y���z��᜿F�0�v��`xy�-=N������-��d�i?N��zG�`�t+C�W�65!�}f	\����K��i5���t锠���nCO��|�eN�)Y��X�cYp��d������1ƞ����]���oO���@B�A��5�2n���߂�D9���N�N��4��x?g�mBp@)IRqGR��W�-�1veJ��b�K���{�L���+�lo���ê�8�AGڇ��� �uQ�oO�T�e�0�M�=���s��3ʅ�Բ�@/��ʾv�f�e����Hb��9\ ��� �TNBL'��SN��U�*�T,Y#� _��H5�Q��`�wX�W����j茞��l�!��O2o�����	�u��!�P#���Fʳ�[�&��%L
��@7Ǫ<4�*,D���c^Ȉ2"��9�S�)���F�����c+��B��F��>K���IǬF�̺��ķ�]��Sc_�A\�ڏ��N	����*2�cH(���9�W@��oa�]V��9S@��}�(�g��W^�2���%@v��!�;�˱#�����n�#i�Ti)-��B��I��f�8�|o:RخK�烳��\�Ӛ9Y�]�_6/��),�J�g�X�r��R��A�>[Rڻ^���׆��YE��q�#t��a_��ѩcՖQV�kX�/&�ؕ %� �gg?�x��/��"P`%Əɍ\�Fuj�����w&mx�.��	��r7�=�^�� �a�'A�	���e)G�'�U^`8q!-ѫ%���r'P�^���Uo%(����b7�쌱X%bc�e��v�}lIi�yP>;�f>҉#�4ѵ�i�mj]���/#-p�I*��F��-���ܧ����J��
�zԼ�����H��BB�km�d����"G��Q]���ZlE[6]�p��[ե�3ess����ӄ"[�L�,��)�
Ro98��yW]�vސ-����g$����s�c]%J'�&t�iAG�A��Lf־���6sm�����>�B���ZDP��5�|
G������&�����I���&n���D]��.�K�}]���KK#qXkɰ���@��<?�ͩߠ�lH���M58AU�n�S��|l�9�4S��S�d�Pw�Ĵ�F7Z5�Y�Z"�%X��o�7�tH93�#��s��W:W� :˰���M�V-�4� ��n�L�OC:N�&&��<�`�&U��#�����S[����Y#��S��/��)�k���G�\�*���o�tR������7�u'�%fq�E�7�z]�fP�,{��e�����5�]`>��� ',�m^��4��Cb� p�%6Ty��?� (:�0ā'�lk�̲AUP��{��l�����Y_�5^���Op�o�-�@|6��5������{��sp�E��`h��lM���]s�O^��[��-Sa>�P��4�`�!�;�(��|V�-��4�I
g<'�k�ۡ
mL���_+ʀ��S�����	#}XM\qp��Z �;��>ˡ�d���j���13�x��|������������S|�l��]о̀R�(�ۮ쁀g�/��?!V='P/���NM��*���qۚO�g���	�հ�?�%�a���ѢżZӖ/�-Rc��,��PC���7"�-��L�B�D��+%\Ѻ3�7m�Jh{ĺP_]!�����t��������^�0x�
 ���>V�\_����QwNo�(~�3W��
��oH�Ӓ�t��ya�Ny2�:�©�����?d�H�{8���o$��MU�Ķ�˥Q�?`�=���0Y�<���|�,U���=�jc��M�ņ�ؖ�*b��0�-�e^��Q����s/���h8�2�W{*�ևp^Z�P�.��:�n�l�M���A/�*2#(��n����;�Nﰲ� �vK��i����W�'.�����5����mA�L�ڴ'��~�j�Fl�"�I�"{E�M@����G�,r�d�>�q5���ʊ9]�ѹۍ
���ªD�}.*Ԧ^�ܺ��r��zJ6�itUq%����W?���7����@��`vB�Un�5�0M�T�[�94�h7+u��v��Mv[�&��6�g��0V��+�� F�����	7���&���)�Vz�� �f�H�2T�	v�5�Z����0rH�����f��~m��Am@�F��ť4��K��|��~Z��%�J�������L����"��Q]�Z���sgGQoӐ�Of)��6HdX�r���U��.��kۋ��'�����үȂ�I,���Ws�� >��L���e�\:�ݻ b�G�L����-l�XG;I/��Kk�� ���8�I3�-�-/��<7��D	oK8�j��=u�r"���5��3�8rG�?��R(��Sz`�^��@�D�����7�W�ڡ[�e����Wx�$P,嬠VF05p}~��|�͜e?��v/yӐ�E#�)�IV�?)�+��D�ؑ��W6�w��c��4E��*Gv�!�����ψ@o�z�`���s��K( #�M�W��۸͚L���/-M��Ht*����j2͑��	��jF�/�1��6(Ss�/g���V%��([�3��S��p����ը/w��nD'�s�z�����-��g[�U�69�*�Mŗ�FT�p��ە�v�6�S�I�I��[���P-W��>����*��y�s��D���GR^��������D{��a/��=|C��u�8�¯f�=��.6�O}k�Hӣ����B�`M"������H����yWO�c����]/�+�f2�]^��<B���#�u�j�hc2�%�ɠ�lR|�'�P@���أ)�����vKi|�F�������/}壥O�Ec�us(�cL�f��ۮ�Jq���K��S�kNKp9*�X}&�����$�Q���܏�%K����[��8�8aکy����(�� �W4a!�g��t5��fy��榄��G�s�Dް����b@� ��S¿c����~�A]x��8�}= �`�
����Or�����I�\�D�7�*�AAN�{�oI�y��:X3�l�}<u��&ӽ���)�� u�P]Z(|�47�t��t�/>�t��y���J�xy�UX'���x�t%��d� ������Joo��?���(ֶFa�"p��u&��D>=���@�o�k^�s�V�j`�������&ϸb�m�O����|֫=���~r|����i���4���Z�o��=����pȀ!�>U�K�7�naZj��q���S6յ+���3m���'�����7�h^���!�X$��6���<����_��bƶ�m�;���������t�ƏE+��n�? ����H�����9�ͼ��*�!=�7�c�$� ��AP�b�7�ʴ�q���A��eq���>�3���ur�.~���Hl_��vK�Ŋ}����;:�a��D���7|���.�>��2�gԀ�>�r��V
��G0j35��bm7�n�?L�B��g����|��ڗ��r�{cܞx���kI�7!U:��j'�n�>H��o��̛�>o^��� /&��>�{i��]�����y	Li��~�1�d�)�c��\۝�r������I���V�*+�|����#&%�=����ٓ��T�n�|/���WRf>P����_T&��6� i �ncT�^�<���"M�Uw�qB�R�^s~�S�|��V��Jx�B3�@I�� �꜎!i������i��=>�1��s������ϪJ[$�����81�lP�I?�x� �4��ḧӱ>sܑ�r����h�-ʥ?F�݄$P63�#8+�rޫ�a���h�s�����HS��Z��a�'`���JU�6�'ss;+��֬��F�u��>�<2X�������t���0� 0bE�������B*��/��/��dS��n��}�0)��GNDye�C�-tH�o�ze}�,[r�Nj R�&���=[�,k�p(��m�"�Q�"F��>G8��ďސO�L�L�Ȁxk�?������B>�"��$�w�m�A���4iˢ-�AB-��A1(�8f˂�h������\2a���U`�](�l��oW��l�t?=�cS	��P���a�h|c� �r$��a�α�$|^6b� �O����b��'Ź�vQ���r�����rw��aҺ�~��y��L�A;'aL�G�E�w�`#9�b���q�5��vk�r��� �D�-)4��E����a�x\'	P�a�YQ�Iq����'������p2�n����iv���ی��5b���RV��sѓz{�ۧ��-�l\Q��DAқ��ۿ:]>q�	����GC��jב���-h��=���n�"����v�˞a���N`��U%�rMJ����X���f}ݶ�PHs�܁F���ɐV�8��o��;8,��=�G���'��\���ᯬd����dy���gݼ�`j�rC)H+ �jCSD5�6ؚǫ�ݦb�������gB��,�3@1���^D��s�R����{����R�5�������z���k����oR6��^0��qa��'H��Gڳ	�$�Zf�]�P�?'�M��*�ŋ�����
�(�jم�����^��˿؂2��Q4�O����BË0�9XsR�!ܬ(����!���6��:��VN�g����Q�i����(.J�}�����	�q%�v��v� ����М�yز��"ދ�db0ĳ-�R!�p}v'� �}�1�TI�̀;�kn���L���es�����\��Ym��+JPP<ma��"���]�t޺o\D��%R��-��͢uXL�ž���վ9�8|�/\�/>���Z��Mw4�=Ĕ��36�r�����>���C�z	!��kz�=8/z�gbqh/g� �5=CK�s��	�>�!*Ks�:�_#� ��ڔR��q��K�|ZC{pk�R�7\��Z�'����)�����`�#ä����T��pw'��&�� ���L��Rv72u���i�\iYŞJ�ILI�谞8�N����n9�TgL�l��PJ|?0�b�����J���Op��=��Y��^��'<���n`�Ӝ�]��C��cZ�W��Ť�=�%��i�)���7/|�O�6J5��$�/w%�*��y��!��oy��TSGѫ��ob�YۻE���W!T�Q�_z���
8�je*��Te/���Smk@E\U�i�4'�n2�4�H�P�����U=sT�?���7R;��\3��亅�e����"`0�@��#kf��پ�VRXѐV�>k#����lz�_;��r;�y��o��Z��zܱZ�^�Ene��['�V����ǑI+�c{����+}Ua*b�D��n�I��i���d\�T�q�����8�mhۜ�l��H�W�i2I�R����A54�=��:��PӑK7�1�ފy:�!���x���І��>F�j+�g���;4Y���0�t������8�B���#�.�qy�iCxl�w�������B}�ޚ9��Ll��Y_�.L(+Hw&nW������ϠW�
�>P��Z���V��~�`wAu���󠫥s
k��o68�#��C6,��ߋ�U�ʌQ�х���zBy@�8Aa�UX�DA�SEK�l����l��zOM5zXc"U�0^�l:�v���Snj}���$4x
!W�!�R��{�y�/eN5��F/J���7�!�8��%��W(C��~0O�.�2h �������c�Y��RyB����a%�j�ҡS�ƃ|٤�}OFM�"��-�|���?�j/�6��+���\��!���nyH	Sm�B�E����He�"@�����R��wcs�PK��x"�Ѹ���LSQ��U�x�-Z����,"�x�@�������� �&��q�#�4˳Sp- �Lt� m0Ź���m�z��T����/w�ʖD�eJ�+p�Pr����F$e͵�� L�PSG�$���˹�HUmKb�nRR���&��ZJ^ߪ��ހ��s�b�Б��TƆ���m,��,w�u�QjSe��z-���]��M �̢�k�*����#eV�Q~H��b>�2��{ ��A{�m"j�i}Y}��0b�vi@�d:w��>F�ZE^�kj����]�.L���$O���	�(w�8[�7B�:�g����権�a��EZ+��'���7�c�.� Hc.>B�Ν��=|9/j���cg2y�{�Kb��>��p�k�F��hs��i{Ia�(d��C�X3Z/[�G��Ҕ�l�ذ�r)Y׸�)�w�u�f�m�97�S}o�eM�Lzݏ��y����ޝ2��R�PE��u(&@��G���昱��	��|d�ٗ��j����B��f���R�6`?��3�Lܹb��N�2n�=����e*×�V��SXG��x�θp�"�oH_�$t��C�xe8�$�\��;�ȑ�:�x�H��D_�S3�h�
!a�<&�kV���7���%�M���Fp�=e$�w5\��16���Ы�����x�b�5�_�\�z��崅�L;K�8���'�Clq����?\É��*��G^�mfl��Q������8Ҁ��������
���f����N��a8�&���R5����-)[H��P�)�24�Ch�I�N3BCt�S���&d*���j쬚����s�<kP�ؙ6{o��E�~$�
���[Ee�ד��S'VͲ�(�q���K�,q[r� ��"ݐon8�H��C��W�@���Nx��J䅅,���r��9��׷l��1�����!=�Z�)�p��� ����(��8�>F��Uzc ����_a-1���k��qZ�jz܁J�9 �o�ы�"�������F��|���P/��T�d���;}x���`���q4T�M��ڡ�P�`�����]'�D�r x�w�|&��w&�S��B����#x�E���"n��a1u��&�m1����_��]8q�*�<7������g�j�8���}�9[�4��"�ј���i�kK���|nly��Ǧ��*ܡV\��2r�ʖ�g�{�)�L�`Y9��h%x�u�Ly��T�Gv|y;����mc���֭1O��>����q�0��b��3��\�R$����$B��Nm��譓 �>�����i|_�0�&�Ӛ�"�7�<95-U�M��a��t<��䚱hX�S������Z?�`�8�YT�����;�Sg��/]]�lR�Ұ���9ǋ��H�KՕ7�v�p�Wt.��_!����t�-K��������TD��.�
y��$7B[;��IF9���������y�L=j�B\���F]��mI�}P%�^zZ<�� ����WP�|6�0�w�?��pf-~�8��N�o�>�����c����Qo���?Rp&T����Tgt�8\��`n搜
r��l�BXFܱ"���B��~�p�iT�]ĸ����#�s���g;��\�Z��^�h�ў\�/�iT�!T�� �F�韁g��>�7P� G�si���a�֓3H����g�\���0���ɻ�%�[�Z�ݯ�}Н�${
�$�[l�H�6s���4��_k؂D@ZU��j�ډQ���ԕ��l_<�c�鋖��)!3�3,KZ������n�wݵW1�� K5q��ʶ��'x>��
�y��d����vg��� ��;'GL�N�V�Qah,�j�R��s1���/�B��a������}��́���±}�牵aXAC�U�|<�zk�)RV 9Ԅ��+�}C�A!Gw0p-����	4h2�$i煺�{�g!�B����+nӰV�؛*7M�O��Q��F�)_�����,���,�;+�aV�ת���z��5�n !*�j=�I��xGY�5�����Ee�����eZ\�����b203gp��;�,� �<�_� TO~���֬T���(zV��Q���uܢ{���t�y�D�>tp�ޒ��ϗu�L�$\�B�Y:D�O-5��\,~�~>��e���<�$�x�~��
*�z��-�J[�s<h�n�kk`���2ǀ|����U��Fg��6�B�c}�jD�wa�Y0�f";�ĦM&w`K��ޏyߘFP��<�Kh��/�އ�}��G��D��sɺ��(�ks�n��o�-�7.������=El�8����!�P׻��ԉ�0F1l�ƨC�Ė�1�!���,���ϘI�g[�>)���a��}��!p�}j�-��M݅����g;�e����9y���u�ƊY �=5E�W�c�k�)o�w�L��63��k��mXj�t�}�a%n�+�
��ց0K�zi�7� o�V����>��!�᠉X[r�S��E@�c����,Vk
���rG����A��i�Bcn"Ϫ5i��W .���b 7ɲ}y�;%��æ^�3%�������\sD�HXM�;Z��hd~v�C~>���O�_���������>F{)�9/���>�ޅE��,{��!l�H����腣���+}�����G��5�DKt��8\a�w�9iD����J���A�(/�^jɼ�a�>���8�l$<tO܋c�1���!K�H���~�\��Ay[�l�� S��]�jo�ߓ�Nh~@*���)�Qh˛5S,�s��F��
�K
b�t��灛X:��4W%j�į����~���vFܼk
;��`C�+h^`�;po�0*N_�-��w����1�љ�"zk�{)���n&X]�	�r������/�ЁN�<Ah]{���K�z[oa	_L����qfc:ciG&�<P�՜�s��tO�Z�5Oj{S�@���ŵݬ�WF��� ���v�vs�	��Ivhi �rX�9��پ�iB�P����brֈ�E��4!��2��'�5�����0��P�1�	���n����H"ee -衱"��2u�T�L��{$�A�>�P�唬F���j�
�e/&<���ĥ׈xr�E��נ�|��%W><0I<
kNӛO��/H�T�8e#e��I_h�r����Z��ab#�!�q�O��(��`{�g�)=�ۦ�3i|�
�^~�Hr�����e)������ϱHr�QY��F�[��o 
f'��OP��PC���� �F�л�T$�����X\�.4�V�������l6�s�eS\ݶ�Ʀ�PWԼDP�uT^;��\߻�K�������x�t��F<���mW��6�:\��\�?2��<�B�fgG��I��~�R8�|� i�:�iƊ�r]�E��uÙ�Q����۾;Z��F�0g}��g��;�W�>�"�<*��r�
N^��s>�� ZKD>��`��B�+C��Q:t}�ר����hKr���L��$���M��>�X����c����_�%~j���)��(�z�./�"!�[Ng )�ʒJEqS#�Q=�On�yi� �x��~�K<i���6� �%�x�&J�C]�|�sd�����i=^4���]������v����~sO�"�����$g����Ѹ�`a^z@��xQAmܮd�[L0�[����k�'����G�HO���੿`���!�$��
z����hjc<Mf!��}�
��/�g;�^L��k��0~��;���E}��($��mR)���w>��Aky��MWԎf�5�J�@,Fs��+�Q�^0;��w�Xԗ4D��w1�y�m_�kqK9Oi�j�t��s�L#U��^����v���.L��i��j���}�?U�~�_�� ����g�Ĕ���9��ʝ��k �w��Ϟ����Q��{`N+�|C��Ul���'��?��_���<쟺0�	��?TY�O�塸�"�Ʀj�z��$4q��h�8:܋)�.:���?e�.�R�n�䶕RN�:���7�T���0�:�B�y�T������ɁT�3[�,fw{��X���IOjz.+�9�����*��>,A�s>�t䩊�?�D�IYy��4�z񾏴=Ux|��ɍ���
��4=�O5	��M�Z4z��~�CzX�rUo��c���T�a���k^��_�v�|z�@�y&O1@�W���� _Z��4�Xne#���8�sγ�/,�ũ	��u`��S���BP"�R��,�X��K*Wо�N�Rƾ�h�<������z�#��Z'���5�X�ˀ_��i����Ik�da��C/�����s�Hgot��Ao9�
]��4)L���L�
���եl����LFK�'9�]�{��;��}#��a��{�,�����+�ޡW�ʬ��t�yۏ���0��O�3�6/`X���s�b6~[}BR���UA��/<�P�ٗYT��Gb�c��5eW�蔸j���(��	:�J*��F�-g�����%m{ņO��.�<��/؂��.�����a���Yb@����Y`<���V���0�z�Rm���O�ٙ����Xh��Y� �%	<[�I@2�.;���'RNn�n�c�}Y�[��&vխ��.(Q���;�K��?�P���b6��u��4	�'�;��4���X�~���Bϟc�D)m��d�Z���m������Ak;�ALM�GẌ�J�C��Cє����m���r_91��IӦZ��%Y�&�hI,�^�Y���]���]W��H/�]5�'sJ�J@�>�	�V��$D�/�@�+��k�pqk�XoS�	ۺ���%�'?�������z!�P�M㥌6[*��eؒ��+������R�D&�E*�[5�2�s���}�Qx�d\�Q�c�y6{r|�ɼ�Z�B]�م���:jYKy�毬*��C���r��ZY��t\N��ӏe��K�q�,6�ժ���)7���g�/ _�r�܆��9눺ʊb"�OG��}vE�Hy�>v�o�{��ZH����ۭ�4�e�����	��w�u�ɋ�מ ���'�35k�mGu�K{[?Ķ��:w.]�;[�����!�[V1�&�����|!-���Gi��wx�\ �Q܆��]A�v��ڜ�&R��kO��^�v����+{%W��<��u�ECOh�vi-�Ȣ/M�FM��:�� �<��S;GM:�H*:h઀gy�g�Tn���&Ay&?jnNl0��9�@��q�>���H��s~�ֱ�O������� ��ʖI;��0��Kif6g�T$�(m�
�	g'f6��Hgn��8c�'���d��,L��dvL6����g"�_�B��+U�h�HV�)����`S/A�K�h,e�_3[�<��ڒƚy�cUv�r�	$�!ۘ�o�	�(�/5fi6$^3ܔ:1�2�q�HW #��۹�cg��o.�2Y��딅h�s�����+�����3�kiDm���v�k ���P8t�5�hih	N<����{zb�=P���>����*w��A�����J�������Ǎ!��7����e��Q���r�KA�0�Q&�d� �4�������J�`�e,�ҖY��nq�d\��mgDz:�V'6�55(/�(0��ӓ9���$N��8%�_�ೊ"'?d�u�]zC�y8����c���]��3����u����u���,�lX�s^����RƑ���V�:Ґ���#��� ��M2ڌ������H�rr e�kX�B��R�[��
7�I{r��n���C�Z�{��-q�l���&\�E6��6���E�ߋ?�B�����:�3������*��	+�BL��<�0ٞ�@��+L� �^d����I��h9�Ha�uxjhE�3�l^��״���љ~2�h.h%�=
3WW��s~���hynn.�����.��]��za#z�K]��(�A�z��;�!)��r�_��r��-�;l�5� �.jhqi4��� <>I����w�r��^J�H9��j����/qQ�}�%��!��6�1�b��-H~S�R�r�'�J�L�A�5�>�1��u�L�K6��	�̈NQ�9�A�[:\.�u":��Fu!��rl��5��0 tD`*�-�yN5�+�LX8�*vf���g���"
 D��e���=H��I~[l�O�_z�H����ʌ�*X�x��4��ϰ���I�Ժϫ��3�8�'�Tp��3jH�����ۡ�&��!�>���P��t�-�p4Hv�� Sg�%O{����[�k2VxF�n:^�����h���3��aYxb�^��2
g*>K����*~�$���/�QaC�I�]+���]�:6 �҉?�܃U����#�ےN��/;uc�8�˕��yU���e�f��s���T������x���+�(�(���@��M ��.�	��hJ�p��Z,�6���r/[��T?�4>�( n8�0I ��6�JOq�g
����ϻ3-�x������4Zٱ��ޭ� �tT{��,���
����hw�����L�	�]��@�n�	�!	S���<�q��zc�^>~?F�=���0!���6:��s�v��pƉb�?�Z����p�d��ME��׏�����ɗ���������,��j/��ZD��$�0��$ָm|2yf.�X�1��>�T	�Ì�7Y�n%�����yӗ=�|<�:o{�6�"+��W�> D�Mq���zT[g��՝ǎ��|�<)�p��Z���s>�|��u�E�9;q/W��1j�0��M56G��U2f���N4���C�?��B�҈�-<��w
@���?@��nK��HDߞC��y+ ��0L��z��j��㹗}y��/ӣ`h��
�]I���7҂��%̤5U����>
�Fg��KP�`-��q5s'�Ք���F�xPF�sYG��A_��YB��o���ܿ�`�ݺ{�Q5�.�J���h]�RL^��V�r������Cw"j���O
�=/�7�vso���]��x�̏�|��r$��^�� ͧd�,%���C�n�p],��`W�Q�5W��騛���_GFt��NE��1TRʛ+j&�ż.�HD0�l��S����
ǋec��[u�?��8m_���?ܠ?�a��1 �S�2O(ұ-N���M��rO��1�sսԈ��d�Ґ��lY9�?k���s���]|�*y�
�Fi�\p���ik��T}�9Ң��u��v���N��=�&b��'=�])>��L�5�?D3�h9HE��;=�	�G~�٦���m
9��
��z����J��K3��=a?R��X5]����"R���k�8^F�h�.`����7�G���6 �Ci���F6����#�%D|C�bb1m����[Po�vO�(�����7;��]0d���0y��C~�K��]zJJI5K,�*�A'@�}���o��Ra��X|�AJ^�����
K�ٔS�3C���l*�
/o��5����5BY�3N�o-(W�P�>�nl�D�'���>#8Ф��P<!ڨ�bDl謂u��}�->������ܬH
+�>u������ݳ�ZC��9�)4�Y�'���mu�a�b���Ҋes�ƃ��mG#O�ހ�A�칱h73��6Gu:�63e��|���QP^w);Ipm?�}Jt��;|����Y�ꈮ  o�����m�}0x�r+<BIy(���tr�O���ry�uʼL6�f���^�2U�pLfV��|4�ab#���!C �m�Z�U���ML��(���Rts�>�xzL��P�W�%��'�&�A�!ƹ#��!,�J��>Z\Vl=���M��q�Ѓj#�Q�Wuc+�M���󍄘����r����֘<n�{�vIb�ZFLK~ŠA;r0u��(w���qE^m�+����DL�J�kl�7���}�XM�Z�F�F��c��$h�2�\�ߞj��))�a�&Z�4����v�Юr�f_L�m��U3�S�ұ ��y-�������#�@�OX�x��֝��^=I}<v��,�P��M��|��QD�,-��+<{F/���-��)�����E�1i�
����*�����Kyås�XH�=��d$x.�����:��c�oY;R��\�k�A9H3g��5�eq�^z*����[=$1p�֌lK�[8�n��󍐾C[����ƨ}��Zv�m-������.<��K��w��]�SV��Cţ�=���b�����p��yܒ�kG�w'^��`�^�0��/�x� 0�ا24�)��P�dK?�c�.�͔e�~�/���2��o���]�G�:�p���ps�N�&:�9��\�@�^��6�O�U��l��z��7��r�P@�����[N.9Јm���3,A���\,��ըS��#�������#K��ix����IOyK4"̱
X̋ɞ�C���/U�W�q�q�Cd�X���N����JO��$��wJ5_�E7�'brޔ�&ji�>�g�db�@�1�%��w���q��v���}Ӊ�*s�ix蓧	�$���e��7a�@`TK!2��2���WA�9c	�$�O�3��kM��c����r�J�z�m�3����-�a���r�4m�=��,R륡����4!?.�Cjp�{�c�r�q�����o��銠��"��7�����kb]��r82�~��d��D���#S��2�,�'%�y�����BLb�_�B���h��Ӌ��(���B�-��hz�D��)Z�~I���A�0(B�H?�h�≟0M���38&��*8G�hKM��ʤ�^����"/��φ�/���˾(�N���'���H����� �uJw+i[s�p�r�"�M�-��؁D�8y˰�P��4φla�aj0ګ85�]���H��JGJ'�@�W���|jyh��`2T���!U�C*5ͱ8���vZ�uVC�L4-+�$Nw8Z����	���`�����/���TWEי#l�Q�E��M��nv��2��[�-�!���k�B0\넑��ʁ��f��p~'�~��dC]�-gB�<{��:G�Ba�,j��]�kE�1��4�䴭Oف���2g�u�-��߮(M�ŗm�/w=Ә:���vLBw�$0$m�d�Q�;O��4���-��׌��h۲fZ���vg�ͱ���(�w������j�����=TGOЏZ�"���`Q����
�f�ǵ�k[n�8w7Q��ABZ����<S>�V��sG�6H�0�������6.G>��@���SD�o�(�7�a��_���������ξ4R�-?���x�0%z)��0�c q�N�+g2%���ϥD*��&e�\�;-hL@��r�?��鼹 P޶�[ ț�k��>ҳU�atv�y�e_2&8(�^}�5����B*r�����6��iw���(K=M�눴a!N4���X֌Vh�~͚#�e�Q�c>2ׅ�SjT��Kα�l��S]��S�`��,!/��Q�'Q��C����F����A���1<;I���d>kD�F�� ��_�P�����҃v���?-C-s���|�;y(�z�Y��%��$#b[ML��Q�K�Gm�^ɩ��Z�������v`�m	I�}�����-hxEΣ�������s,��2y-���%����#�$��,��sb�TJg& �%,`���w�޸��Gh#-�3'���tE�� ��s��CD�͍��]M=�R|�+x�%�qiߊ���r��.6��� #~ve.�qA�H��rC�C(9`�qG�_�GlLC�v�9�W o%�`�1��#_4ю������&<��р��"��a�q�Ik`?�y���-���o��a?�ܬ|nL*�״�z�^8��[�w��b^t�;��$�Q3o�<�0sPqn� ӱ�0��T��&��׍�}�SI�
s�5�i�iƽ���@��H��Ao�ǟ���~�ʹ�0t뫃�hP'=��-n��9GQL���H��.RY��"�j,�����)��,0[�2Ȗ�L!�f��uIS�F3f��m�H�Lv���1kL�[)8F�\s8�e�ށFe ��W�:�-��z�$X��: U�E<"��������S�H?n!����f>�sL
�f�F�H��{��Qr`&���|�a��U��P�qx�:ߨs��"�s���Y-z(����"Am��A*�)?ׅH� m����z�ʢ��`����b3>�9C���h��d[̡FQv�d�S~��G�����7�X~�+|Jwc���F?M.�EGY��[��а�s���80��l��Fj�	?X���� -x?k�{ۤЏ�f�5�|��t� ���{��)W&Ww��R���Ud7	���>��z��|�E�x�Q�8�����7�/�L*�L.�L���e���J?=i�Ԏ�~�QO���R!lC���U�c�";7��g��q�DoK����!1��=��⿮G�G5*�*6����� X��D�;�㑑��LXE�|��(B������Z�GC���7���L:�7��z�_2�M��=� ����٬�'2�����n��R���Y0*[�iʶ)?���Ҝ��>Q�6����T+	eg,n+Hv�1�V�7D��@�Zz����bO�����U��1���Y*�Z_��bxµ{��&�g��^��h��/��@�-���4q����}݆�L�!�3겾�Ap|]ק� 6�F�C�:�Óö+b��x�I�H�x �IRˑ���_�4>��L���Z'|�҈��NJ��!b�c1h .��A�.!�	��'L5��r �f
jK|\�����L�S[m)!��AZ�^�%f�d+O_]����s�7���n����uD��F�v~{g	����0,�r�b��#˿��al����x	��4.X�,3$3�0Za�@�m�>g�K�����>dg�����~�x*u��F���V`D¼�O�����1P�d�.,�]|,�/����y��[to���w5����y6��q:ϋ���o� �����P�b���d����!g	hm����}r�g�m�л��J�GF��2�iC/�;B�"2T<6�'LC�]���t�@��z=/��*�>���0�P
o�͜��tB{��xP)n�����ӔG�Ĥ�nt2�{��L�$t�1f(�O��RA���^�EQٗ�%�� �v+���"��+3�k7���,/*�(��Lo	���+]�շ^T[�����bZ��!�*��F�j��BP`x=�����!����05�u ��o6w��d�2Pn#� ��_��'���A��� +��Aƾ:�Oھ�.�z���*-�L�KA	�6��E�����ޟ\7��Qڵ5?}��{��uy疗]#u�P��FX�(}ʧ��� ����Kpn����e���gW��N�g)����	��*p^J��AMK��-J��=w��Bb?Z�2��>	8u�(�i|�1�Թ$��xrH����ޮߺ
)�xOQ���\mU�HYxDg�ZK;k9ط��1�Ĳ����e��B��KȢ��;�����_�w)]S[�)�YYC^&�u��s)�o��;��
��f������%Y9=�4��J��˂i��PI�}���̕�y1�uk�￷�9�w���5c8��&������-Aް�N
JtW�0�9��;"�BK��3g��v�IC7��3��#��Թ��Á�Y�/�b���ɣ����=�z��Aa')Z�vlܦ�K�}Bhxef%�ͷ1���F�`�c��u�ʢ:��!�Df!�]�Ժ�es���s[Τ�'�O��Py�`��`}Sa.{�)����Cw��BF�8
<-zs��GeiC�/۰�J.�.rMId�}�9� ����$ �7��k��s�z�5�����U�w#R"�����y9�V=�!�ȓYO ��}0P����C}��絮��{�nHP(�RT��w�O�d��͉�b�S�`A�x)gH��[���(6N]����ϰ��s
���~��5(�^��6}�c��g���f��*8wˋ_�׊ɶ Q?�� `�٤P��W�Ve����]��Nk�F�E��l��܀�bf,�1s���~�����kʂ�y,)���篊rw����xPW8�洰\\�D)0���LFpp�:h�&Y�h�2p������8U�<rh�4p��ж��j2��sz[��9���D�|֗0��������S�����?엛��#�})x��T�T���<����^�#B�5�H�U�l�E�j�R��!h+��rt
��t���]4o�V`<v
��w|6��*���`Ħ�}s+E4׎L�:y�����wDא�ݜ�51^�!&VD�3�_�0��P��VPvr���@js��\��b��]�U�$m_�.�	9��NL�n�u���&�S����p���#�N��罴r�R�zy�JAq�RU~�1��4P��~<�����O!�̵ ���T�g�Ǘ�����~r�p*N;B�9LG`�>�m�aF�F��a֨�Y����]w��������7q��|�n4Yr����Y1�rI��DLF��[fM>.}�9=1XkV*���=�u���T*o`Ġrܱ?�Qs�u���ɤ�����=Sx�S���5�k�$:����@�c�YOD�gFEiU���R1ϟ���:s97 �MA�_�vK���;�+J9x��S��g�>|tـC�%�ow�]��Pc�U��������������ye��?h��?�6=+��e� ���q쁎�����+b��fZwh�sp)W��!q��ڞe�VON�����G��դYsl�����V��z6둵8��3C������WR2�����+Pj��X��6e��FN� ͇G�)����y�:x�+���p_���S�/�o	W�i{�5��9�m�����;�Yæ��z�:o��J�~�(g(��(E\����,��<`�析H�c��^��.sR��Ƹ�;��Li"�
�;1u��lM�0_/�	p�4oK@pUC�
&��g��YU}���;u� -�B֍��]d�
>A
��F�\T��~��.�����D)�B{C���l�	�L��9��̕+r���v�e��z����~sq �Iԛ��e:��1)M@U,m �������'���IC�a�c����&�m6eC�,��%�+�����z��ץ�mMe��;SY.�6��j�VB��P��^.y:s˒Q	�绊��MY��������z v��N�3��Q�C���]i�M��ĺ����7
�պ]�S[�]���l `���R�M($zI��6���%uWR84.���^�f�o�r�����`�Ҟ��v^���7��K����q��X-��ky �62�}�`?�1�=��T�`������a�2�f�(RuK�"r&l��P=��nۜ�����T�'��L]T��kf;۔$�C�z�-�*��p�+{%��#[ܯ?y��hX<��L��q� DR�n^چ��_gɐk�KsB�lbZW�\炦#]'�t�+����0˯;u7� ĺ2-��E��iϽ����2��	�-͍�x� Ñ�:P�z���
��pE^�_=� ���fZ>)y�qF??���q�Q̙���$o���B3F9b_r�!�h�Ȼ�^ޏy{�,�yiH�vS�~�_=am�r�U�Sa���ǔG�<3�A�!�ux]��"�|�;���:ti�Z�����-�^_q4�h�PiP��ZU�%��L�_ڮizؕ/��� �`���1�i��\�oXYWu�?��5�?�$?������1ݘ�����'@��XUD)����ڟ�d��(�T�%��K�`�IAHi�鳂�dͬ����@�^�[��'��
Eo0`åW���U�C���jJ�g�Z7���(R�x>-�@�V�P{�V5�����F�&�4�+�)��p@���Y�1�va_4���c���;���v��}W!�6C>9��t^��ˁ��,1����=�[+!����5�5$��:K�J��+M�T�ߐ�����[��y�F�T���Z}ʢ�݁-Y�&ka���U��]� �@ ��U��(Jp�pTyP�C|��e�>���*E31&�A���/�^�&�{Z)�.�f(uFB�ʹ{����f[�S�2���1�mT��?�ջ�����D�;
'L�4-Gul�F`Z3e��"�b��R4�1n-Eƪ���:F��$��ܠ�����bk���ȕ��J��~-w�/l{f���w�U9O0e��6ЃRԹ:��h�N��O�h���Y�	����J%���G�u��s����#�騿_��bIW�pٻ���s5N��sQ�*��.�� �I���T���x�<`���@6���UPSw�Co_&�6ݪ�%{�ӓ~M��BL��';F��p8�\��g3|=��$u��֖�*��G~�[� �wOT
���~XPP����mʩ�K{���t�b��{��B疑X0���t��*&>{|�}�+��VP��xD��i��ȦLm��[�	<K��
X{��~|�m��).0�fg�B[w��F��i��덶D��a��I����A`��G�������1Tdr�5�hd��O��[�[����󟐹�;\���Kg�E�(9V�����<�����a��N&��8x;����>���,�+�w�����l���B����.�����&&l��F�����ʞ�:+��ߖ�.����O��SFL��@�i(&����5B��@���FrʜR�W��\���(w�r2�$T��v��~SA��hYpP�,��?pga����W|�����t��� u&%咄��)�ৣ���F)�_�*e�#�c%�m�j���%""����~=)BQ��`�U��s�(&�� $R��[z�� {j��4�Hn�쾛Х���8����}�^��C�C�_�`e����' ��b P��Ȓ�<�^쁮@{gM�}rp9�r�(�������P����Pp��?� `�CZ��� _՗^E��K�{"����mM�4]��_:#K�A.�ʲ�Z՛#�PO��e�9j��
��Hh�Uꩲ��h�d���^E��{Q�`�g�s�}���ـږd{���lٙxx�=���*���p�h�~!!@(��?%.��9�xpY$0��ˮ>z���}�'�˧��zEr_Q�u#���'߶7�6�Hc�n�!F��{�)h�+w��n�Z�0�%gW^k�\���xw~x�sM��ê= G`�
:��D���Y���d���Y�������4pLɞA���K�wy��^�t^f�#�,ʆ�A�m��s�ϋ)�&�Up���^:��ݏ�����B
^�Zw_H�}����pwB��p.��g)&��pi��n4.��y��,�N 'nN!�t(:Ћt:��]3��n�H��t�_����	WH� a"��+��p�u���(��F�M�|V�F0D������A��^�Z^Kn��P}�m>�U8`oʒͩ`0�m�6W�XI��tt>U�y��J��! zt��i��DBˠ���#�����e��\y�9��-�2�_R`�*�{����R-	(�oI�N�x�EA�A^]59�g0��T���z�e���d�qq���8"@zJz�)�����д�b�W?s�� !�=�~��	" 
m��|���{N��E�1K���cL�A�Mn@�$AدI@j"z�~9��;{�殚)���܊�T\R�q`a@Q~$C��!98/\�S�ѓ�v�vvE�.�����7��^��H��nIya�V�BZ"�\�+ԝ����L�rڮ?!�s	���br��~%�P=寒����#"2�]:C����̉������\�ə�$$��Ǻ���q��iT���,�O��8��Z�M��mp)��s�  �������4�B; D~ͺ-x�f������?F�,2j��M�1������U-@[[���o=��يu�����ſ�A���D��k��
򆏫��/�*V��U�9�)����6�zo\����n�(��7��m���)��4�H�Q��D�N��O"@���Y���v�*�s�)�/��Us����ƐJ�r��߰��]>NF��\};�a	�b���d+��7hkW��w���Y�����Ekdĩ�:5���&y�@��n�NG�!�����0q��&���=���ds�H�i�8����3��mg����N������W�}(Z��C�4�Ib8HL���C�LIP�Ο$��{	�=^���`ϯ��-Q8�������'������������Js��BjT.��#�TW(�:��c�}��1� 8��;���6�@���zCm+<ӓ���y�4���6�}��&ԃ�T�$*�����#*g]_ޛ�:#�Zg3W����"���۪W��E�����j`�D�.}��E��9��"�����Ui�h(Hp��/��#y��D����`��Є9[����K������~;Ӌ���Bcd9����?,�����ބ���d:��/|�|dV���bzS�=v�B{���2�z�*���H���K��?���\���!�� �;�PV��+��{3P䕺y�&2il|1~��\��9�\W1���_�HkU2�����.��[�r N���u���E�{�b�[]wH�$j������;fETD���&b���0�3nl���q���Ԥ�2(�-|�'�[[}���L���˴�`����@�:�U+4z�A
lg�q��B����b_�|w���ы�Lx�K߽�mH�@�[P��/���Ǻ)&�R-��Ҙ	7m@����~��yp�wdC��A47��S)0_�T�֌v73��R3%����>���h�Y�}V�Lq�y<!���4�OI�7�!썚6/�?���wB%��`���]�j��:M�6�3�+�>���E$�����Y)1ӟ���Ɖ�R�0�5��ϩ�|�bwȕ?�b��h)u!�yԏ꫶[��M����Cy\��G߼>ߦk�����ėWe�O{&X7c7�4"	��t_[`��1�t_h�t�u �?�}���bJ����c!4������8$�ce!�-ނ�x�F���o����6<� �/b?�D�v������x7]�%KW���ƥP~ji\��1������mt�*��J5�2a��|�2�Y�Ǣ����q�2���
,lC�L�I�	�l�;;x��;�n`�Np%�N�TR�u��{?+?{�o~(�이a��2p���m�=�	������y0�4)װ�ִ�hD'!�/ &������� ^Ӎ������C���y[�����x�'D*����E_�:��9��œ��yGV�k����,�T��ʏٹi�D����80�)�:�B�7{��3�5�-q�E)F;�	�(�Ӕ�:�+*h�%v(Y#p�� ��3�Yg�I�l��2iȽ����t��Ћ9��%�}�c�5V6�����A�K(;�j��-�C��O�L )��l'w@�ĪP��b���S]}���5���f2�3+��OBƒ�_��q2��/N(��5ŝ*�Ψ\��s~���E:H���3�]�3_��,���i�ޣfQ�6���I�-.�!��ś�\=4 �Y$}��+����Bq!�������,�n}�6<��e�o`ד�
{��d'X�;�2�ׁ��������4��Hp����̡�QQ��g�
��x��V�|� �k�q�4d6}���/yK����b-^6�& 7k�1�����n��Y�`��cBrX��ja_���oc���FX�F���Ҙ�x*pu]KG|�����_�N��:=lb�R���3��|oh3;�5{��xQa�\�N"��/?����gŘ�4`Ujz7;T@��קz;��ʚ���%��Ҏ�4Z�S���5dJ|�����)�m�j�T�@�Gx��2$e��<2�t����G�'{F�ü�Α�U�z{�����#�{m�C�yMVr�61�><�^��L^M4������	�"2pv`��)h0��y+�������a��y���m��@����^�=zѡ��h�Y��e>1�9Ћk�߭O${����2�6h���Oq��� N�j3ݵ8*&�Xn�˝@�T�G�T�[} Y�����+��"�~Z�bA�p�����>����x��f�ۑϤG]R���0�Q>��e�NJT�/
�ֵ��'�zT�gP���� xǁw��p�#��c�([�Y�qY��H��GE,�11�j��������7�"�jx�*@ȪA�J�l_�
�/�	݄ᚯZ͡�r�#޾��`��o�� �me+��K�k��>��~�	E�pf�Ze��	[R�%��L@M���k�B�l�⏮��p�hh+�����+ZV~O�V��4��ޠB{��P�)}Gi�sE�@�g�KV�qv��Q�1]X�az]����&��׬D�Ʉ;��n�8�q�O�+k3@z���4�e�p��0��b�Ƙdv�6Gk���b��s��v�똈��l�0�`��]F�W����'�:F*c�[' +>�r�����L��^X@vK$��1� �U_T�6���,MP�v`lp�k�����gBA��v�1�&HP<!��� ��CK3��N$�E���faHP���2���6oO}���"\4]����{g�gbQ%d�ɣ�%�J���u�h;%x�8�5�sx��,G�bkD�,Oj��̒���SS���#�KxӵE�!,�R��D�a@j4��r�D
i��M�4=6�N�[����׽�8)�oH�Q�����b��4B�.��Lw��ٓKUO�r"oW�0c����vi2��2����`9��gL`dԚӏO(u��� ������ �aC�@&�&~��Y���1Q�Q�q�`ȝ��˖�n��R���2eS��R��
;�#�xM��Op'����:e��1�訵Vݠ؟���z}���J�9�$�ˣdOo��@t%�'��pPH�G�r ���b������T7�h�ڒ�/R:-_Jq=7��o�|�Ԍ�G�G����`�[\��������z�dQ�2i�E�6�r07��G�N����B�ZDʶ�=�9 _��V�V�.a��z�K�QF���O<5��#�^ 3%�ȝ07�$d�ڷ�����V����p����*�e�����%If>2����jw�l�K\tE%qx�2l��"�-v	��M�׫i���9�Z�˱�m���2K$����4����C㥮TK�lu���g��LV�����u�#Ŋ�袟���tQ�f���h5�-���0�q���.��<U˂�+K<{~�p�qGF��l��Ǫ�g���Wev�|@�¯���#BSe4u1�!m*��M���=Y�[Ք���6`����5C"?T`��F4"^�RO��27V�9Z�]g���.���I<h��T0�3o��Ks�.;;��,��y(Ϣ�^=Y���ȟ(�*�St��nwֺ�X��|2jQ1��XoK�Z>�T�+�5� =\4�$���<�u������{�o~�g�:�=�U~t_`���ހ�?���{ݮ�\_x�K��;Rd�_pKB�����9�Y2$�_�3RL~�e`�M�8��hg*h�B��Q�n�7J�Z_��% }��d
X2_<�ei�0���Ê�����<eS���!�4=˔�<���\�,�M$�>ڃ���T=�b2fv�#^���}\�#�n��E���\�jH,�~��ؽ�P���w��UA����v�,�M�!9�\J���
7ɱ8ԓVl�-�gQ����Y0J�VW]v��| �+���]��^�8�w;����+��n�R0��Ǳ]߅n5R��=����[�
�:�-S+~ϓK���z{d�;����AP����c9g5e��ǉ �@��R���fTɚ��5���E��ȁ�l�	S^8�_<W�2��QZ����b�(O�M����R��|
�`�����+z?���>��Qi�L�N=�Y2S��&uֹ
�%��{E�hF>�l�X�Ki��R�=W|�'�q��q�&ަ������*�����pߨb'����I���~U�HK&Oss���,����Fy�?�yB�i�
Q�w�"��!s��}�{�-�s�1FpR1���hP��mQvdת\%V�q!��E��t-{r�N� ᘿ@3�$Og0S�_��B�--8p�t�sh��ԙ��($���ICI���ͫ�Zz�aq�N��|�����0�@�V�X��p	TԆ�̇�׬��j���j����PoR�n �=zC�����4��1BG��N$�� ���X��
"0*7�:%b��6��)@o8���4��\� ��:�nmT��w�X]��|�5H�JY�S.�=M���W/��>�C�����E��L���YcQ60�����u꧌���j;��A<{Wm?�H"~ˠɮ1�]#�L���5�3lbN R��q((>�MF�XH��K����s-Cqj��J"�i\�̩z�Y�����j�ΐ-�Ԁ+�����˼og��$u`�:�:��!�I�x��O;L��3J�� D���*>���d�ӕ"~a�qhep���+�<zj�v�5"}�m� �FÄ�T�UEӖ��4G���ЗR��;���o��p�o߸ou *�y�°�� ⵩��'���Ķ����O��j,�CPx��4�l��՜"�I�3�s�m��E��&*�&��ڞ�n�%�����������)��uw�:1�o���x|�|�ͥN��9��2��r�8�@���X�Xg/��[?/�D�WY�T@
3��Q��[��Do��*&UP�Jc��0e�+�~7)s�) �����<co�ے\�ڷ� �X�
r.?��+�a�[,p��T/��cz��}��6m�S�sCR���̭�ӣ����[�*��Z��kکk���tR>���[��A.*��@S�6:�8bK�-��]�0�Ht)�iU?~��+2��te`��-j"�KT��i+W���i
3�}s�跜T_���C���OB��x�IBv���ٞ��M�X]j"�X�ׯ{#�Q���|�:"�AK���:��D�q�f��{e�}��~6��l:��SDCdu������"�g��O�ʘ�H�]�!w�\���3���.�ǃ��B<����;��[�N��\`�c�1�o������w�)0��9D��Lj3�>�	���<�'O|�o7�;[j�C� ��5��D��Q]�r[?���mm��md�]�K%XK����TKf6���/�3s�l�kp�.��b�4\�͹�q[m�{xp�C�Z�P]��5MW�{˗g����7Բ�T����Iԝ��M�����M!e@@1 �T��^��(�
���Q�[��ʹu���o��h�lh��Q��8��C�H��z$�dKQ�߭n���\2���~'O2wO�3 ��ǘ;v��_Pb6Q~��n5>O�:"?�9s�༾�aZ�C��,�ԱA��X���	���o�S��H�<<����X����SkS�C/Eau����(�J�&k���=���Y�xZfx?u|(��ޗu���ԗƗT�:(j)�_r��O�g}�/�����%����}��,�2M�p�����H4ܫ�iM\r-S�'�a1`�Iv�\k����)�U��%���� 4��G
��Gr#�M1�)�oT��RNRG��;��q^E!e�aXi_��rF�w2���^���v���U1���J��k�� %��.KF���&�e��b�u�#K6X)3S�wL��9�!����,�wd��&�׳fP۞%m42 �{�����zǲ�nj�c�i V�9���q��~v0lc`�A�C�eA����!b+����!�e/�zS���m�֝Q���fE{�#?@�wF^�%��[��n��W�p�����(����x�:M��s����QF�V���ٯ�x�s�ꦑ !*��/���Ԭ���9�j���WVKD���#쮢�ʒ�(+X͖��k �����e����|�bE�]��i޼�],�ۛz�8��BD޿���\B/GWY�����H�ܭI��z�ŏ��8'�.�A��f�OҘI��P,���Ş���:�m>�;;��u����a��s�T8��t��?�)5�:W�edfǶh���KL^���S��G�}�3�����v��06�'L�
荗�k��}�����u�Oc ߰��*47i��k�c��5��E���N��WBEĐ��a������l�"��|����Q��M%0hV�&�-]�dxr�L�Q=��.D��ycCR�&P:�]��!����Js�4�w�q�')i�P�2��PO����T;�	��Ǘ��M�q����=Ţ��CD?��b������PQFS/>�ضؕ���SUߏ��2����v�	�B0*f�?vU��Y&Tgz�wxP�e �b�1V�1 �ms�\����,6^��	��`%����3;3���7t�v��3
��WY	O�9��p�Zhn̴�m�,��nVm����;�����x��6�(D2�޾U��j���~)\�	��^ߴG�zX:��D5��j�Ld+I"�(��TPD����曏���(����[��M32vĥ{�ے2B��)��W9��䕱GرE-�H�x���PF.k!�Gi�{8���?\A҅N�e�ݐ�����8�-Ǎ�}	xf D-��籓��A!\�ݿ�4��e����\ʮl~�Ԙ���ͥhG���~�eU�9=�z�K�9���M�f���	|�%_�X*����E�_Z�y���.�.�z���-�$�7����X��D��9r,O�zU{/m}��'�6}S,�H���I ��΀yTEB)�cBP���җ���R��������Sr�C���TQ�K���1�����"c��a7wgO��ND+���h��VX"�mqg8k$���{�СX��">$��,
���nʒ��;��Rזdw]
���#L�f�	F�*�E�	rj�8I���N��2�l���0�C��(����2y�h��@��O��6ZF\h�+��2���k4�%u7�R� $v��m�w!�	c����M�>���B�%�gu�����	a����ɋL��{�Ć�ϰb��m�-Q<����M6;�� �����DU�L����/���T�)���G}���-�CM^��R�SeS��|�� ��6zZ�����z�xN۲&������r�n�ќT.aq�v\���y�Q2�cD��m����c�!�?< �u����O�w��	��<�߈|}�`N���]�R8�M��C���sJ�j��F~H���9���C�s!\�	�߯��0\*��Nh�`����/�8���&=��=�8��¿r8�2���Yv%�j֭�2:�
���1TBKg�3ؑ6q<���������A��"�����H�Y5��7�]�0F�%�L��,;�BI����dG��=����;�Y���zyHҿB��=�]��n�̧/�V��5
y��h4үG`I��}Ջs�Rw�1�I-]�����j�n$!�A7I%�HS�iԍ���L��B��������u�~]��l�م:'���~�̝͆���̓�́=U`T�.����ɔ�W���3��b���y$=�D����'���A���`��X��u�4|�jw1}����}2��z�T�h�y-]̫�k¯�Q���֧p$�����<; ��B���e	n��<'d�'��J$�VǄdC����R�%F�ϫ�-����LV�md�Z�۪%��4����-�#/���%�I�,��4Ąk�]p?��,��;Mb�m����Q��B|d�}�RT�T�g���ެ�y�\M��.��a3|T?�c�j"	6B���X�A�w",�A�*��t�!(Aݍ�_,�Ԙ\�UA1{��%�q���S-6��0&��	�^�þk��`�B��]�҈�O�apւ��,� �A�@̅">!�8t���	(�-�6����xOX{ňW�f�������N#�l��q��Rq�|_.:���SB4kiu}�M]1w���|�����TJ��c���!,�����s�^ۜ��Hi|\T}����X{��}�|Z��2��@�d��u� �j�����pTD�u�q���fE�yqw*?.�� ��yjzӋWhƕ��S��~Z����d-�v��5;K,��xe��n�Z��<�����-fHG�*�fS�M��o??w&z!a�)�aY�E�|^��U�����&=D˦;�+���G(0��ec����X_��]A废����GS.J� �k;����nFq�j�IB��A ��e�{1Y����cZOg7m���*�gp��xvQ�=��\����&7�]�H��>b�Ui��� �8���caE�rn�T��H��V���T�ȗI-��E�լ5-�h��I�l/etƁ}^v�6"�Q.��
ފy�i}z�����B2B�Ua�����9k�	^#r �|���zi�H��@��h�

�Ok��Rб�YC|4�kÝ�Q9��q�^��s�d~�}s����_�ִ��ާ�)"��?oxWt���ĸ�qp�2HT�~ңl�i��Ϙa�a~2O�o��UG���;2JeǤ�i	<rIv��s����l����ԅ����M��������*B�u�Y����;J�C�"�vT�C$Z�O��Q\�f��Ü�R���<Z�ۈ�hCƋ�2�Me?�v��N��bb�[#��l�����c<5�,��e�M	��+�b�.�O�_�uY�-\�����䲘��ޡ�����om%�갅�ʹ��uZQR�3�I>��%�C��_~;��%����B�=-27S�+�0Dnޮ�/�
зP�ɯ>�wXaM �g��۶��K�P&*�:%X���J���vᢩA���ʶ�A����Lf�E-�ĵs37�ޒ��k	%�zǅ6��j:I�'��2��'�w��k TNd)���G�<�\J�W:���ր�Y9G*n�	4N,���:)�a4F��.��C�l[��%_�v0=B�2�hа)T�������g<Q٦U"}��qy��HG���i�0pް�JڥFn��k<[�ܨ2��D���`S���D<>���̄�S�����"��C105�l��k�M=������>{;4γ�� e�0����ŃKf�+ù��1>+?'�p���� ���g��:��-'�n+��=_ˤ��1�ՠ]�u}T N����0��<i�H<c��xn�0rP���������>�]��3�o���Y�I�&�D�~�t�Y� Wg��K��<Sw����,��|i�ZRu@�$�p�C�[X�=���|R,`�C�� �A�YH���Gc��s'eH�A��)E���R��t*��I�.�����,P�ɟ�d��������4�dH�{w]?���� 昃�0�	3ǔl�m� N%0ٗ&�F �@.ɛ��ږ�#%5Kω+ʤ��{�d�p��y���	�q���$�uc&G����"nF��.���uw+�A��iWǞ�-��Md�F[��[��\v�a�b���������E������wz�#�S��9r�|���b��� �L��U��%���ԣ�+�Hv���drbԞn�tuU'�<-i.8,�_	pc��j?�p ����cR�*}7�т@;�oT��DSL��r��DA녩AFEw��<W:�ck��z4��U�������f����/U���<3�����3i ��n��n(���~Y��X[Jf��_Q�����5&��������q"��ꂀOeG�Aß̜��a3.~"�E��Z�7v����cK]W���k�'�
qO^�������u�@m+b�%�J�(�>i���E���F6���Y��3�i�M��.�ٰ]"m�c�\	����J�d�p�e�ϘD�#b��ݵ���׍���?S����esB��-�[��Em��qP���~�yqU<��R����1ς���O�D�� �Z^�gb!s���aV\�؎Uϫ
�O�����dx��O𔄖��Έ�Y!�a�Z �z_�=�":�Ņv�#!�C�?V�U���;6u��ߞ�>�����ҟ�M
/����I����i�^���ed�H>b�Cn,r������r������-P�s���13 �́����A����5#���w�f1�7T��!�	�`q��r�`��>Z��B:�r���M���c�T����i�}�5�E{�~?���h�lp��oAỞ3�&�MM;aa�h��b�6�+�}K�f��L����A�`_�L/@���K��W�L/Q�>̾����3;|�^)8�|o\�U�Ŭ��'��f��	y��	x�$M�d�	��@��<���̰X
�b����ϫ*���PKN�U��UH��R]å㧡o���Y�c��V/g#��Wj�L>G�i�n}�`�m���I~I�.Z�-diO��_��f�YhfB�寥��	�i��zArC�Ku�T}{�<��a������E<�������^i|�]};�5�ynv�����
�}�DN+>�4P���ΰ�����>%�O�rU;�eC�i�ʢ
�o�6��3Ŝ$ ;���)���S��x�d�K�뜐Y��7ϕL�Q���Hy�?D�����6�\��߀o���k�j@jѠ�ɸz���Q����T^��6�K��_ֆr��7U�<��[!-�)˖����Im]ǂޔS��X��R�H�)j� ܠ��j���t�(Q(��g8�3�U���.͓���m���B���F��D8/�Sd'�s��kn�����i�{=q��g��\]����텗a�R+�G���B�N�@yB������MDI�^�5~�D��Qp�+b�lL��s�5Nl��Lギ��vٯ~B�å�Vp��g�=M����K�[:�����sO��I2��ֻY�K����n��<�8�y{��:�|�Z5.=7G�k��G�N�AOc��/�-�e&��o廃c��F��(�{W;���
FK~C���Q]��3�Q�`�R���J��B��2�\˱��`�4p eY���p)�}���}� >���$3&�N���f7�nf�M2�I�MM�k�)Q�͟L���ƛ%��X�W[Xc<_6���kփ0�@�8�aa8����B|H~�@��x���H��Ο�D�l{��#g5�?Gw��h�Y�4Ǖ��* ��.yO&�!���P9��5{<#oc1�7N_�'�8
��ߎt����b���zQ�=��\�<l}z�� Ƃ�m#�6oqn��HC!�1� J��`\�DI2>��}�z�V��ᛈ�g��}�]w~��К-x��խ����XH"G�B-�E[���3�=m}��u�{�p�~}&�[V�"����u�B��Z�8�?�Ν���'ψ'\Yp�u�%27I����W�����W�1��^Ӿ��n�xu�sk�N������"�)���s�~��@��L�f�㲟}�qB�����[5�MU�8��c؁�A�?�Г�G�����`�'�f��&��s_�|��U �������<�.�a�Ƨ�R�>ِK���D�yMf+��ԯ���$�$�Qi�tUK�(\8�z��Xy�}L�����R]�ق�e-ַF7�Hb,]L�R��ŕ�NB�7U�J fj���5�,��9|K~E˩<�s��F��c^�h���-||�����(�tf&b�a������^�s���=�^�*���9�٠�TV�I(M�s>�N*A�}F�fӊZo�:�OE���R�{�Q!��wZ@Qu��^�ڳh�;;�`Q�AQm�8RJRْu�V?��a����`���X�X�y1_6E4�PRՖ.����Í��KNR^���b\��VA
��g���(�!���`��"S�oKE�Np��w���Y�b��VS�4��u� �\�@#�ÈuZ�x^eR�8���d��[5����^�s��s/��;�4�v��3��j%ԒD��Ś6_Q�M���#�TZ��M������k�ly�x��^��aI��gي��1�������00�����ݲ�)�|�Wv���.nk��?��J,^�rS/_��1�T^�&�c5&-�����å璎8z%i�!`V��g0��-�\�\�Z�YH�0B6���L�~�8���X�gj�R��jh�`��5\�u����HY�x�߇��g����K)�T(�8�����x@6�\|0p�ֳ'fW(��i�u�s,�t��^L�4�Q��<�w�S}ou����D�Y����9�/`U��b֫%��TN�+�Mb|��-�u9x�����ܙGL�ݮ�G�u�ͱ<!�>y�a:��L��޷cdšB��\��(���c|��.w-H;y%�mz�����d��ғ�Y�5�F�x*���#������ś�;�r¯ZȪY��@{��\!蝨'I��S
-��3�_Z�_Ǧ�z�R���&�D�����S1����a=zt9i$����|�
+b��k�4���]�e�q����j&�Us_.��Hb�Ra�&��bx)�J���/�%y<y;R7�tW}M������!jn4�H��p�8<&��ǰ��dp�E���_gX�o��َ��|�+�{�T��_>�Ͻo�F
��Ok3��P���
u�p.e�=`�H��w~[L��$��Ip�۝��N)G#H����,:,U�����JAI �s�h��^�s��΅H������ʹ�+q�'kPޘqd�,X!�{\f�ݑC�O����bw���+���k�;iC����L��J˜�����s�Uߢ9�XN�w��7�s1�
h���Y�\��Qf$3���6��=�.�l��e\> ��r��#ɗ��Ω�%�$<���6�b?�{d�V�Yt�
�Z�:3b����ޖ�jq�R�򮓴���p-���w8���됒,k҉
$��\���� ���ў\�y؏��1Gg���^���w���<H],�[���D]v-�� Ա�������R�?��&�O��Kq�)a7�t0v���s�%�y�A9�3�m>��Ӊhl��V�2��θ�j��� 8gK(4����u�EA��b^�t׌,q��|ˠ���m���"�X�C�6��⼏��sx�nfP����ݙ������#yu��'�H�.�nڶ�B��-^8����t�1�LJ�O���@�2�;��K����7;�<��"0�����5����MU�����#�2�[wA�3-&��p+떮=�"T�fv81�l���Z�����F�O�\�?'a�Y��x�ٲ�-�j\W���u�B�u|������3��YA30_~s�fu��L��$1�ɔ�ڽs��Ƒ��p�ɶ��a0�W3C
��D��7�x?����ˀ�w�c׳�>лE0\�"�{�e������(�%���Q/f̹`r���ëE�I�2��.��QZ��U%YX�VsaͦRc��b��&�t�&�>R��%~�FŚ[�rhr��X�?�I�k��r>i�X��@>�f��e�A.���O�����<'L��5vUt�vC�0&zI���k�_�P�>�HU�����Z
�M�"['"���������71-�M�=�@��K��L{e�x�G�	 �ٷæً�Rc�h�WgAz$y�E��A���JL�{"m���νe)���N��
�JYK��?�\�^cs�{��H��Rw�r&oz�~��30��u��c�󁦬�m��Lp����֕�u�AS$	pTĵ�q���z�C&��j��<ҿkZ�2�Iz'��l�f�_qC�+�h�z����ě���l�.+�ǉ+����YT2	�@�<w�uiDC��b(����\q3p1O�I��eO��#v��S�ܕ]�~����6b���-1鬪Gl"��W���UuP,���ܩ��G����}t�G8X������"J�af�̜��U}�ϡ2�&tQ_,q�t�@b[<�vX�J�=��p=�7Q�sy��k�K�BT+�o+�O^��#�w\'H�{�g#�s9�"-#�T��wa�0���\�,���|��|�#P觧c��u־�=��9	qHn]�OW�INq@����%JT�z)�'�H��	H�+T����cޠ��mG}q/������w�0�I:#CQ������{o��gɤ;���xd\=�뻙�x��wXsA"��-�V�w�����:����pji�svxjE������t�cYطI��X�j�K�I�������mӰ~W4_�x�R"�W��l�=EǢ(�P.\
�D����;�Ȥ������}%f%�����f֮6���G���)a��6AGT�\����� .@�p!�`�5�z+3	\�m�,�!TQ��me@LU��|Q�����t�Q�~�]X�S�TN����	ۼ��7Tj������C��#m�P�E����u�#��d2c�,��	�k��%eһ��]wsŜ⡩���ɢkuVUaMJ<�[�!��!��5���y��:b�H�b)%M���+hb֔�R �G��x5�"��m���\cP��;ߝ ��M�׾�{4d}��"�{{����0?��l�_噡��4�����������V?�ַ�[x6.a��xC�P��dޛ%q��}��$��Z.���\��+B}|RZ�7(er{��&�V�j�����w�J�iQ�IKN8w��8Q������@�W�]w���%&:Ǒ������R^n��rn�gL�:y"�����;4|C��̗�"Q͹s�I77M�y��⧉�g�Z�]�i��E�s�|U� �)���O����)7�X�,�I�Q�L��t ��w�r���BK�������-0u�Vz�"�ԓi崴�{��r���hTGK�xT��c��H���=w?Vc�L��{���3�AW��ӄ�Nf,'�t 娘zp�UqVb0���B�p1 �[>=N�n�FI(��OX�q��/��s$�x.� �͛�"�	0�	��HRJCϝ١�ąp���(Da���c&��m��׸��W&¬ /���W�ן���CD�j�@�d%X�腜 S��ꮊ'乲G�8R?vU�����z�u�C�'OӰ3�%o8�C�K�0���WK�u��`G��3������sj0�E9��~����&[�g�M��̥�W��Z-�+O���O-sG񛓲6rН[��,��Wb���gy��0�޽���)���N���!J��R2-�`�[��t���������P�?!�F�JK�m9�oi·�ףԞxcLf���3�*x0��V9t�TM��h�)le'���Nt�l����Ŕ`�7*����RҍJ�p6E��n#!�릞��S�c��n\a��RP�����,�j!jR������GQ3S�۰���o�$m�MI��%2A�4:`�-�[��v�^ڡo���S|����*� u��m� ���4��`'Q�VŲ�u^Ա��#c���uƼ:e��R�����v����!�/�e���=�xj���bh��|2J�q-7"����ng�Ad�F_͊�$��j?����u���`�K/wk-���H�=����!~��E�{�,�|����Tdd�j�k�|eF�Q_���<y@6�Ti]l��7r_��br�~��;9������Լ;��TY�"�<1P'��ʳ���CXB�P7Ɏ�hd����2G�=]w��ڒ�RT��p���ި��ŨQ��)L�}h���0/q��.�g2��������eX�M�/P���h��� �4|*_iT+��Z|�ʖ�`hk6�����;S<�/#}��V %U��'T�*�Ꮟ�u���m^�~�z]�E�%U�v���	8������"�;�QSn�ؐ29�\~�^'2��L���f�YV�	o�؛n��|��·�~���-<�!vന�w+B��b�ڝ�]�5z�VHv�*�r��U�y�&��^�W��Ň�ԝ���-	i��0�����i3��gռr`:����	���P+ �/��H�t����Ūt����#�k}KT1ywj�h(�~�8���p���ׇ�T
�a�6�:��Z�n�zɭY="D�9�~�������$]��}-ђ~\��̤|�qz�X<У�ZR>��S@�C��1�ZN\��ϑ�a�B%v0�*�:`��q�$땰�δ�<:�9��ar�wg�:�H�]�,��d6eJ�"�bK�	a��y�\��@"s1ty���_�����q�;�˙s��#u�h�#l�l���vX5y�jv�_��K��څ+���s�BLT���&|6�,��i{H+��]��X�����t]Ӻ.7'ߴ%����/�1��Z�~9��_�?���-���x��"��n�����CDƽ�mbK�?{�et	��F��� /��c�"�`{�����8O�6>y��-�#0T��9P|�<�9�,�AfB�"84O� '�u��k��\�7�\S!B�t���,l��4��ݽ�x�e/��HZ nCX7;�m�_=�;���ч�20ʜ!.?XB�|�U,����3sc�2U7Z�ܜ�b�tA�嬛b�emoe|d� )�S����F������D��Nu�M2i�:3K����,¹��H�E��K�=��AT�;Jv�֝�f'������A��i�NWC�)F��D1z��gRE�̡v���:Ӈ8E��#�@�h:	�U����S�������(�u-[P��_��6U��/��ǼI�3�rdsZ�ꔩ �t� 8�3���7خ� \E��/ڥW�g���.���%�d� ��T��ڠ22����������e]tu3��7�2�(h�'�Β��oL�Y�д��(WnxUWeC�V�NZ� ��hH_"K�9<��3��d؁$?�(~M�۰0T;ɋ�G2�����@�:a���m���.1OK��e�KZ: ������xA��D�AH�҄��XqVV��H�������@|�~4�r��s�!�դu*��[0�ypP��<�O����GGDx�x\6��<p�&�.��x���q]͓�C��P�`Z=\���#=�^B8�����>"�|
�b��x��Dx2qޢ��A����8J�wL��K՟�S�6(-P��A�T�H�#��;x��i)1�sz!�*F�~�?��Yx�k?$�-�l����ڹ�^�xg9�x��9tW�W�n�ν��.�ۄA�z�c��:]#a:&���/��%��_O+w��
JJ���s,�ϭ�3Du�OY���3y��r�6�����<�|�9��̫$8�Gr޷�����F��b��% (|d�H�J�{	'\>�(A��_���!j=45�Z���ܨq��mRej�ҔZ�s�>˭C�E�Z��5۽'��3�*DE4;�L\��S?%-,W�9��X� Ul#� 	�'O���	?� y�!>N�I.���c�*�
n{v��8��7[^��)�?j��W_6���L�P�P��GG�X�y�R"������~e�)��>A%:?
!I�= �#��!�!J�:�e1����ui�I�E�NG��ҋ�
7�B���^2��
נX@g��'��P6�5Hu@1��|&�� Ws`�� �r���f���П�Ի�"��W{"[�?�c�.����4�:/c�/]ח-��T�;��?'c���&���7�g�1�쬾fa)2�M:GAm�b��L*a�DHsS�?@Q���^�kKh��T���@�#�SD�~f#���ےg�j]߉{�߮Sf{��.�B$�y+�nq��u����%bCi��*e/�Dz��r�ބJ��k�7R!T��M�+�@�Z3��L[հ
FK[qP�8�a�_����fB#~�eM�s N�r8禴C���	��6���i՗(w@�YZ�ݳ����t���7&�>��^�)9{^�2���cŧ\d���>�Boq���}Ր����pz��K7�`['����L8eb9!��t�c��n�mcYKI6�!�핳>x�e�j��!����wv���i~��� �i�`�yR�ň[���E�a��3�x�������Z�9>0���$價B��Ԙ��}��t�;@C�I�����C�×�j�M����IEb���*c���4Rn̙��U�%HH��F�&��Wt6�>Q��Hm�$@���҉�W.��ZB�w���`�`?sd���Ӓ��6"6����>@7�<�b����N���|��p���"!����� 1&:QTK�7S�A��Qa:�,�!�3��!�_b�T�pֵ<8ĳ(��{	�
�puf�0v}�<ܮNm��ai��m�����~���ͥ]��^�1�,�|~ �H�n�Tڶ
����-1s�W6�a�)�!�����71sh���v�&6J�Xk�,PA/���x�خ���s�"mܼ*��+��=?���%^�U���e=��(���(�7tVT�ljqR:�)dH���gto�(����ގ���Ii��B4��^�8f��9�܃����BRCw���QwL��-�y�ӂQnKF����>��)��SwŰ�f������ƍ@����?L�pG[z���D��8P�j�1�@�R/$;��ZG�j�;Î�L�v�e��<�A4�V��D�C��lCU��`�
H��R�C����C1mɶ�@d�(e�	�t�[>(۲|q�Zg�#���ѽЗ`_�����j��5�_!Ko�@��V��#�ҙ�J���|Lp��F&/fتJ�{�6�)V�"��d#�0?�{�j��T���T�:��,�2Pua��0�����q�s�qE�֠�+ׁ���(���dn�	�}FI�SN�!�:�a<���w�6��E���9쎍��r�/e/�
��$}�w��P)(�oXi���Z��O4���⨧����$`ۛ�sx�%g��6�e	v��m0�`aQ��Y�k�M7|��@��-�ͭH[����2�ޤ״59���X�ѱ�zu��1kUP��a �>N��>��+��ݹ*��DX�!՚҆#�y-�}}�s���D E�G=��pנ�\v�Tt��C��r�}�C��uh�>�D�Ӥ�����үd�������M/���
�6}(���ݚR� �鎻�7A�2'S�6���.�f*�r;\���Q��	�^�ٽn�T��Mվ���(� 'w��2��Q� ��:T���q�oxq5��n"k�&�Z{/�ȟ��KX��wf��2���`P�t=���2�8a��h�ljy�z��u�"����)�V�J6s�}�\��A����["�S>,���cGg�"VX)��7F/+�g��!����ƣ^=�_��2&H4]՝����^8V���Qz<�--�^E��2���4�d�4��s��%�%P��b`:x>O ;�l����ּ��p��}d�����0���n�k)����u^�1�bH($\	(�*Z�a(2sh�d�d��y,8�f�B7,.qc��"Dj����R�?cUm�,U0��+�x���ߌ-J50��ڡ$��c���>�k>5����oWK���wM���ںOMU�K�S�Q���Fi;6A	�1B!ۗ[�ȮB~�Ϫ%� ���i�@��Mq��DV��1K����WS��0"����ȼjL6s?���A�0�n���GM��Ƞ���e�i�Y>µ;>�mV�������ѹN�&�~�g��mw�WfӲ�-�p9r�й��&#�� ��D�	�=.Z�
ƪ��Ȍ������Bk�J����B.�G'����v3M�Zh ����>�{i�x)���7+�uy��
��[!�v9�
�ؓ��2~����cֺ�q�[2�p9U4�}�K���}�P`���Ew���L�����9
��+�S�q9�/ݯj/� }�Yu�9��Oԃ2MK��5 ]���5H4�8[p�ȧ�|��IqQ��8�TnR�q{8d����>���y^w>��"�ȥN�uA�����p���t�� 8RE��`��y�H{�X�S5�ck���ҫg��-�hH6F��7˸��>�M����Wq�g��S�L��K�ֻ�K�3Ns��_�֥�3{�c��;D�l^;���_�$-�Jk�~��޲#�4V��sE̙Ȏ���&�V%�rQ�ս��~I��w7 �N�Uo����d�}A[�`H�d>	��E�P�+7IE�a�e�*����e�K-e�>%[Lj5*�#T�P���_
{��z�%�%�L�o�pՒ@;��ټ�T���=eGS��#��\��4�ozM��̝$e�%{Z���WˌUF��F jZv8Ӓ`�,�w�� �됔6���߲�t�@3�2'd^z�dP(�@i���V\#p%�A��I�t�h៦ќO�vK��ځZؿ��n	bɓ����6�fۗ4�D\����~���xg����R3�E��}�hٟx�̩��3�������9�|%�͐G����2r����Q7��}�YRؖ�C7u ͫuv�l B%�w��x��\�K�ڠ}\�W��=M^e���yE���[��Vm�p�lِ$��c�f�����1�\��ꘄ¯|���VM�d���>%DM�-6����BD*͏Q����H�Ľ˳�G�V�.�_H�����7��+$1���@d��o��� ���y�k �T�L���|!�k���l��PW��mY�^�q+]�Bb��F8���w\p�x�p�&���k����0�bw����ҢJ�ZI�_�rInf>��ucLs&˔e:@e$�Y�c�����J�&���~�*S�6'��΂�H���<���Yڗ�Mox��{��p���C�����B��cb0/O�� .�[:K���f�ǎ5
	��T/��"�l���Y�K�d]MVKY_#�$����ٽ$dZ��z�I��B���H`�Ơ�_]nq2@6?�~�ۓr�����E7��\Q�އ���3a�Q��;I^�e4w�T$���7����$�R����q��GK���o��i8`ۓŃU��"!� �T�������@���x�N����Cq�U>�b/�����0�0X�D�����	ѳ�����+��Ju���it蠚Ryz��H�9r�>�3/p��	��]9A�s�V��EE�Dr��V�6�5e�M[��}�91��Q��t7�4g+�/X.;�es�.bv��(�	�m�ip�l� W�`J+W��ض��WL�L㒛1�Ui��F5)d���-@۟'V�[ѼA���e�wx%���eR�#2��9.�@	.�xt��'N�:��&fLHn1��N)z�-�^���?��ct���P�j[�=����=b�!���1O%M�X��ae�$����)�|���fs��3����رƨ7F����)�����~�r/�wX�IL������	����C��N��_o;��jU��_C��}2�_�Z,ơ!�fTZ�e�h؃2mt��:����ʧ~�RO�����X�3sC��}3��j�rR8p�7�gi�k(�k�������	��q�O��F���(��s�:��'�N�h(pq��q�焧@���R��6J+��4������K�S�)��XNP�V_�	k4������N�<����v���A\t��M�rH$lT2��m9tveJ��N �1�Jm/:+��Ҧ�2��OU�K����y���@rR�(�ڝ9�d������5���DaK��|�2�l��� z9�y[�8�I���lW��@��&��!C���*�ߊPyJ�8��V�d0�x�a�4�qYw�;Q8�|��lGya�]0HqL'-n>g���y=���t���՘}�_P�Gȶ�Ɂ&M۾e�H�:��-3qU�j��و�ߠe�v�(�8H4��^�����)T�dkXc��D{��
�9���8���1Z���>I��rGI�z�S�s��ҾȐ����cX�A�������/�KS��k�Ҫ��n`\��n���D�/gUKP�=I��e� A3ҟ��{d��}e���C��a;�׮LzTI꾵ʠĸ������>����p�|\�`�<�����;n<f�$v.Ogz��.����)W��[u�.c�U����e.�b���N����v��1&�P n@Ӛ9\�<��0tB��ׁX�Fn�x�
�l3��C��)�)ڎ���9oj�»%�4��7f��n6�Y��E�u�k�M'XY��,w��O�D��-��O����C�9h�3���U���Ȃ�ҟ���I��S�<@��'^dSDR�wۦ�&�3�_�k���0[?_��u�5���G95&{��I������s�W�e�~of�P�p�@ay�.���xb$�=pB%๨W����cOX}GN�䬈T�{Zm�-4�Y�8���-�.k������'I�h�D�Y'���]zc�ϔH&;:�/�� f:�y��,i'�N�B{-!2�k �������=����ͯ����U-⏈������E;AqE�D>[%�>��E6��<�,H��ʆ]�=�	v�p��>�ٻL�a�����(e5đ�G��mjߕ~;���hk�ǊX��e���[0.F� �'L�'�_2	��@R�vA�?KynŘ{zYYɍRO1���}6Gi��(+�� �4��oM��7p��OG%#���6��������ᆿ����<D���<R�(��5��.�~=��՜�8u~�����nh縗�!�eUbZB��]=8:��a�&%:� �R7[�X�'�:g�Cqg�p��>Fi���'��@��aL7q7w�_/fx�y/Vu�AR�y��C�<A��=���g��8��8':�C�F�q&�.i�}���|����#��14ӓHR���d�R�,��a�ў�t�S�
#�Eh=P.Xeغ����Շvn.��Ϥy4��m8>j~���=����ąfn1�*7f5���T�h������D�6�u:FC��a��ƻ�\���O�ھʖh ��a�����+�vEW�N�NF��īܕL�sZ:%��@�[�}P�����������5u�:3�� ���hp�C�T�}���A#���� ��#�bu�7� h%�Ø�g[�N��[�0��u��-t?Ș"��D���#l��?���+�%��j����;"�P��8i�U6KZ$>�g�מ9��2���V��<�zX-�6��)3V[͒��絁=�a��!���sqy���à����;���C�<M���~�v�>�G��,0=?�T��iaf�"n�Y�^��k�k�F�L��/p ���>��l�?+��@����~�yj�Z����κ��_��iP���r���h: �ys�=H����Ή��O�vA��	~���{�������%>2�����FMa��9tG�~��wb9�O���s�ۨ@@Ka�����Q�Υ���Q����k
yT%��U��b������Agݖ��v���S��|d`�4�p/B��m*��!CFA��	%��&lSu:9��KHU���6k�\~xه��;4�F�s�M�RNËA:���H���C��ul6d M\u���1�����8���6����z�$�]�&-�3�O����14|��������v�cY�a2�XM�|x����NE"�}��Z�^�&�Z:A��#�S��[���#y�����lz�(�T����$;��><}��.�&,T���*�gb�K���6��S���F��l�7Z��󾊄k��:
�;�L�����s�m5W�K_4�v_��R�s��H!��e�U�򠁺z#�O�Bk�(#�e���4I�.3�!��C�Qa�w��2Z��4�K�ɇ�5�bZ�t� %�"pA�D%�f�}߈/~ĩ.���Y'�au�Z��b���޵i\�!�]	�HV�ၚj��-��E�q��՛�"9FG˰DB���/�SH%��bJKֺ���DѢ�R��]cO�lk�7�_��g(�-�zi�D9%��QSw�ϳ�|ݑ������(�?C	%�[���!��lw��Z=�/����Ӭ���ה'BM�3�m�<v�S�㚨F�zw��/���}	le9�)�� �^R5�e�s��1�jSJ(To����Q�d���Ptw�!��l�Tɓ����v�o���Zx=��M�d?��B9�������lj�,Fp��u4?׻p�!���B�ޑ��x�1_ۘ�ԮFϑ�	;.ƏQ�_޼����%QW+'��������'%B^��q��V���������A�����Db�m�f%Aʂ(>�OvP"{ꉪ{e3Z�$�~�H��Uk�EuCg/a�ı:A��Oy��{��K�K�o�G�\�[��m��,a��n&�V�;��f�t48�	�ۂqA��"s�»е����:�SSR�a�a�=�w��Ҹ���q"7Y����/��wBn���04�ʫ��})E]�.�;�w�A;�E�9ih˄J��g�o{�igQT��F��[Z玵\z*2459������*~��`�!6�s-��3E2��Ç�]��U'�.���Ǹ�E�E&-s�@q?���F(G���[k�?d1�؃�7ǝH�I���z^���*�?�ϟk��l]b�ɿ��U久͌��0T��]Ȗ�Ͽ�� m�Q�w�B���b���I��(���y�t؞E��ڥa���C3�~���3�<WC�E�ǚ�M�[����s�x���q	�m-�^��\t��'7G�@��=��^��C�=������|9�9����"��Zz���ר1�ڕ��FRA8��*���#��
A;�Q������]ը/�_>W�]싐�'��,*����p����'�m�0�8-��a�<�ML��c�����8��Ppz�Z+��ĳ�o��ў� ��Ȏ�!����_\Yy�~�_2�^�DBר_G����x�mt�f�� 
0�� �8��L��"�U�Zb�&9��+���deX��pbS��rz�7��wѾ�Ũ��
;֯�����mV�����ά���=3}7`�,����+����2�8T=�lWx�"3�.�}��+a���u<��70/`ͩ4��v�t��:�%Y��$\�����y;�R5��mP����E�7(�~:�!X��Tzr�4:���|�1E ���TG;oY���y݈W�wt�@)�	ا��[@�#�{��Q}��ɂ��2������w_��*nʇ\lu3B�`�̲�G�ΚCKA&�!P�̤U�c�����٫_�O�$Ci|�[B���Գ�\����H.�;���D�z�_�}��������:�cT��\�/"��ӌ����v�����Ҩ/>yK�/�5�3���|�1���=��<��<+M�wjB��|����M�=`xj#"�m9"]d��L���G���!�0`�Q�S~8�qҥ:,{}˾|�x%���Ms�P������M�/ ��l�϶dk��vfKw�vҼǀ�'v�i�hn:X?�)�_�����{<Jrj�Ȫ� P��.�w-w����q�K��,z�� gc�������_�۫[xH�.��e�k2��L����>E�����4��~?��<k�������+߇�T���Q�F���)�bM������d��F<F���A|�M�b���-�ȗKKv�e݄Q�)�X">.�tعa���!A?@ݍ��E��|ח [�b�r�͵s��x����݈ȭ�^���IP����%w�k�̾g���|_;$\?�ؙ[�!E�`j�e���Zl�9z
�K�ب#�t�b�v��5z���2��tv�R��]^��|�i��?��F ��������k�Z���I��!��!(d�)�W�Ҵ�J�U���J����(�܁.��x��64-��>)���om���u��eg�i���!LL^���y �����v�I�ݱ���\�Nh���<ɴoft|�BS<��Z��2�yu�/�Aj2��%�ɭH��=b}iM�njt����^�I���4�W��j�r�Fu0�ҎdNK�<2E3}������x��(�فc�=��(vqB�r3)�B�ݔ�����eb�)z�&ؔ�A��0���$�F��F('m�њ]Zރi,�҆�*[�b�I�W�\g�����[��l����,���B��6�5p�Uoz�4�Qo�h�#�*𷿝�F���K�m9�����^Y7R��L]�0���͙@	D�pE���Vu�{?��.n4�G�m�0�/����2�2���o�dp<?�JDG�������g����}󨡏��l�ਤ��oܨR{�6_��k�lt�xE�����s�uܷiw���S�=|g�G�L~T	�.6gyh�{��I��7+>�"ot�S�_�'v�h�%R<�.S�}W�by�����I�'��ԩ�Ѥ
VY��e`,���Ұ��k�S���S�|�d��,P��:��<���D?�)��q���g�.	,���|��N����\��o��td�ܱ�~����O�b�9�z��t5�N�F���!�e�d�F�X`���f���hV��f���
Z\�U�*��)q�^�4�m�YGys�'1j�:U)ل�����f�d�k���%_�ŁRvj�n�O�yYя��}_&2g��S���^^�F@�$�)����/�{��~�@�5��orn�BM?�T�5t����'I�`Joݍ4ű���|B	���n�:o��#�Z�����\�m�7&F?�W�;�h�m����j.� �䣯����� JТm��99�q�������w'�d��? /��/W����f��E8�����&�:
��5}v�dJ���i���8C�: �������j���+�0"cR�5b�]5�=8tg��>f-�FH�]��_�XY���C-����c�*�1!g����,��0�%��|�(�I25�*5�Mr�:��c
�v�;F�P*w?0|h#Wf~���.Vj�g<2��y���	��e`� �=,	� 盰��,��o%eqe�R�H1�����\�)�(��|��җ�^���Xl���x�vؔ��{�Fڥ/� u-A�ũ��(��]�m�/#[�Y�e�p�$Q���tL��'J,�xp�"���g����ޠ�������t@eZ�R�NPpnL���"�B�E����	�t)ߢ`�X6��}��w��+<ީ��׫u��Q6�'���0�hsx���6�_��� Q�"qʐ���qF��,�M�;6+7��:�#���&\��-��9xjK=>�A.E�y4�����a�����Q(���8�E�uQ�2[���K�	�t4?6@����Ur�����W��hFR��S���YU����'?L�Qc�=�D�L`�B��{=B�a���ލ�lv�pL!�ZT�xF�Ġc�J&��X �i:�E�4��F�{�?���%�2�ƕk�Cid,����F�����{P�<�����N�w#Ͼ�$Z�O�Z/	}-dA�=����yN�u�X��<��X �[m'q�Ηw�T:���5�6(j���������s�;�� �K���Q��^�A%���ɍ��Ʈ8���\�9^i�i����Jl{*bAv��@���!yM�Lؒ���/]�Rx0����LxT�}�
���o~����"��&�vc�q�	WӔ�eTg�P6q�;� RL����^k�H�#S����C��ЖѦ���yٞn %9�~���\<i��1�����6�}����چ�@bx�7�2�0u�p'7pO4�%j�B�0$�J|4�HHU���I"��"�\�A�j�8kHu�uD�-�i��zڰȬ+�R������� �a��w�2z�@�w��5��O�1Xp�˵�k�i^Тާ�c�+�r|n�	��*)&��d��ˈ��`�A���d�:砘lV��*�W�q"�Kh}c�j�|�6=�b�.�7�s��~,�k/[�3��@���8�xj�B�ܹj* ����,&�&�4��U����IÁ�.vF_�?[��P ���Ɲ1;��ø�naº(�{�u9�&�H���U�il�%�
h;�ĵS�H��
� �����Ȋ�L���0���Z)%t�AyJo���e�}��I���!����=�m�!��3]j�U���3Ұ��l��l���c܉@.Ԙ�'A
b�t�l��oa�#!��#)P���Dv���b}��'Qi��.�}����:���-h�we��7�.ũ�l������ҟ#�+r�{�z��H��E�=CfN�$у�!{�4p����ЄZ/���\P�:U����i+�1_*0�V��䎜�ݽΌ���!�į	�����nMr?�!�$�`*��o �O�G���.�������1|��M �O^YY�R��?���`ܨ/�s���K��!������?��aZ�*t��w± _���{�G�Z��3�B�e��U�S#4��x@��f�-������F{g�9���K��ؓ�[��`�h������3h���ԙ��a�SF������zn���l1�ㅆ�nNmfŀ
w�
f�B�q���v�ˎzmiv�n&'�3C&X`N��WA�y�5@Ѕ�w��� ��q�-+S�bEǍ�Iy3D2l'��٢z}��W`H{��v�:�/��>DWF���I�&0����[���s'u^ּ����F%- �C7~�_f�p��zܰ��pK��/nuS�̺�M	��w���{H0��;��E�FL~��u��2cg��+��
v(�yA��*�x0>,-9hTI�J���(5{���Ppp���/�@r+Yq�E����q[�nW9� �Zc�r�V:���d�|�=Ïd�8'6������/z-�G{+M#�uT�Kޒ�T�S-μ8y�@]�<��cm�4���˜����0����|O��Lc���Ϋ�^]y%��2��j*L����ȓ�K��܈*��(5�gBQڝz#�m���L��#��A���uCngyRȤ]*��S���u\�������}C�4�)A��;��g���?���ַ]N��}ߓOU�ʶR�U���R޶��L���$����X����t��^9]{� Y��c�;�����͙����c5̬m�~�QhM���UT�R����q�N�n��"������m�Ѝ�
}
Yh�/t�<ǶS� MK���c{�#�V+R�IKB	���A���)�[�}�^��WC�U�l'��v�^<�e`��M[�-�t�K�Dq�p���0r�7P$���0�`�g0p�g)��<4mO���x��Ka���I���{O¾�>X�n�M_�h�z���t�4�C=c�Li�^�-�|=�LQ��k����Z��z�U稇)"���AB���U1!8�@�`'��U��HU� ��߶�Ĳ_�_̦�tc���Z�KY_[�%�3�eJ��yv���(�X.���[ D��,u��J��`��QyL�����lf����:�ǯ9��f����Ӏ	}}�y<_�Ou�
���sg�0��-��3��I?m����_qg2�R˵���Dm�ń��mo6]����0j��S���W`ǰ=�ܝE�P����?��rhX�\B��>�H-�'-�dy	v�6��C��^ �B�����e4�Mڭ���Qw;6����^/^����;ڀdY��Z����k�l9��Ҡ�5"͊g�=�Y�ش��2�E��L�}Dxoa��2G�u�@\G���Eo�V�L�7�$��i����P����ǳ����EO����|&�,��J̮���QZ3J���5��:B'��������0e�:^1���x8M��X0���l��K�s$7wx)����A@lYg�Q��a��hb�τE���!��H�&l�7^�#hsj[@��Ɏ�?ߞ�5ot;\�k�D���p�Q���+��Ü�b�Ru(�!�����KV��Ǉ�w���UΈ{):OG�}5@Q�y���J��Г_�r������ӭ �.��l��������c-F>�&��Z��K �xj�2S����w�_Қ҃�uȩP.xB��C�y8�������6��a@bf�"t�y���=��4Cl/,������:8Ke�������zf�Ջ�������7V^M�.x~��(�(�9��e��v'$,�]�چ�yX{-�����Jᬑ!��L�oA���Ӛ�l�p�c`(�JL4h)�nY���S�_@Ў	���}�Ahb5�EA�����8��F�=@�E2,��Y�m�L����<���� �t;����͎-���Y}T��2mIl�:o���ȣ�k�Ɣ0��i���9��[B2�I�w�D�s��(���9e�;���"�"1NR��$�n;L�>��	Z=�y�ҋ���4�5��H<��^��>(��黜�.�\aAv~��5����g�]/!9�ӑt��'XunR� >��5d�۔ȔV�*�M�-��;�{������JF�����&�iG�?-Ѫ�&��Ǯ�~b5�嫁��v����IA8�{G5�/��ocd4�/a�{��,�Z:rK�1�Gٴ���L�鈇q�ϳhtz�E>]�qݡ�y��D%dSE�K�D������xW��`��Fo�_��(�$.�O�y��V!D��@�Bwd* cZ<z�^}�A����eq��(�3�s�bN��������|���<i��?����:�æKo$.�h��m;�~o���ЏT�v��Ć�ݍ/3���*ή�JK�z5����N��8${=�^�}+�_�۱&Y@���-��p�s��*�vkXYN�VΝiW��L�/.#/��ڱzZ���ى&ԴNJ�je=�7Du�9O0Z�ރ>՝A��o���2�$�L	�6(�C-K\�����T�5<�i;�`�����9B���q��pѐ�cA��;��_Dӥ�ҡ��h���/|�hD���Gq���:�% ��"��a�v�w�th)��M�:y/s^C+HE�����7 a����W'H$O?��!{��Hd�I�a]?�����ݦ���_�@4�"k�G�
�d4H�t��z�V��B?��>Q�� S�5������(r��Ñup?�atPS�󄝨�c��n�O
�{�v4��>�ɵC��Z���a?���!Ib�[��l_>t��K�t\ʖ��?�\�QZ&���^�
"�4"�x��h�KK��v�I�����0z������r�jo^���:Ȓ0�el���s;�`�p}�����*�����i[�<%���/�����`0�ҷ��o���Aa�����1#	�������u��4��O�q��jp�(k
	|��uT��Ps#5�r��S����o�˄;�ZO�z�˵�ĳ���Se�4���S�٧�[|�BPJ�c'0��6�`j<�(�c+p���O�J��qk� H�u���.�?�n�	$B��kh��b�Y�5>
B�.v�`csܛ�n�"�Eơ��C�XS�?�W���v��K#S����U�x����6e�;q;�����ebg���{�8؍��+�խ�Yo��?����U��%�)�u��iy�����y�,L5�V�E�&7�T[����_�\m�a�L�{O2+�/Mo�b�5�6$���I��X����ڤᚔZ?�	L)�қH��1����|c�Wu�ٷ�|���(ü�&H��rX�(6^��m5ˣ��<T��R����W� 4���mq�� �=�¤k�E��,�p:�b~�(�-��w���n}xR %҂H�#��7�F��� ԅ������[AcU��\��@:"���±�-��c�R�6-�H$�nW �;�]��c=�KI��Y���7��9��q�v���(�4ZMo�Rp˱��{;Ey�-/�#��z���p�B#�@&�yM%KIh	#�H�O�^1gD���*p��g�S�*M��o;�W��;T��H���G��=IP$L�"�n� ��h/Y��r�?�q���LkpFO�@�׮%�4X���F0��9��P�V鍶eY�V��gc34��f�[ׂv�vx�		�>����&��N��)�x��&���d�e������ǘP�����a�y�G�(S��9V�n6l�\w�z�>퀹^�K(�-����n�V��O���R���b7���GB"��E��7�:Vn��8/^�[����:ަ~ �)q�j������\�eʜ���#�'�-qǆ��u��.mW�����ڳ�?��J|(^,�j���� �	���!WwRi�2CtW]E��n���|��^�~���>u��v�{�g�RD\�r����7��"��9�u=��pxxM��8jb(��	�f�V-�q��+Zh+��m܏Y���7EɷpZ�����m��vw�����7˽�Fʯ㵆�z��KY귏�h���v����P^����HK͟P�V;z p�wy����U,RG��5�n�M�c����T�)��o���e�t���+��r ��K=���fTe�EI�򙉍kܟ����;��ל}�t�%M�$�f@�8�;�3�.��=�ӛ��=���f�m�d��T����B��S�U-��eg`������'	�ɥl��Ώ1T)V] ��9Y
ބ-o<�${T��{'}?��$�GԻ�0���:��o���K�ݡ������'��PaK�S�k�wtTWTh�V�_��"礚�edI��<��y�G��T;�!���4I7��$[�iFa��H�F�-V<�֔o��n<�j�v~7Iyp�! -�ϥ��p��!�15�x���_V��.� ��<A8Fk.}�OQ��Xn����� ��a���o#A"��e؎L�=���D&����$r~�k��&�z�AC�{�"�Ll_�U�@7=P�~��&�w��gDi;����P�J��F��}�p��n�-h���5Ii}a��ڝ��t�݋�C_bӐ��=���+x@W�������L���a����&^[������r�yh�D���a����'���&�A�+d�QڛkF_.��/���S�e��mf�����,�aZ-w�����m���PC�u�a[R�4����b,I/t�UL�)�b$�y=�7)�9�9#n���G�q�:���^����"t���3~��"��sKm��OM����z�_�g:Sֺ&7�^��{��������to4W�1�0q�B8�Y��J���yh���v��iL,���E.���"2.".6�H'lQ철�jtf�ey�[��f�g��e">���_e�����[�����3�H��M�r��Kt���_�u&�O��b��5�E�G�n�v��:D���@���^�����޷tn�aۀM�p7�5�*�R}Mܱ�P��R��M�BB8MJL�j�#A�x���FR�R�NK1q8n�h]�ΔR�Vz���Z��:���/:�S�3�JpX@�3d��֋�O�n|��oڿ�z�bψ�oǦ>g�j�k�b4��hP���<2�X�>��c�8�׋����5�"2��T�v�����<wg\�j�L���5R�C�w��ب���UƱӸ�K�
���Ѕ���f��yQ��'�)�("�T��	�z=�5�  �L��"c�^O�>^psV�P*�Ͳt�˰
TK'�:��Ȣ�(�2<Bn,�/7��2�t�F #Z�]�Bgb����]���G�-�] bZ#?t��İ�i���r���y��]��BD� ���`�J�G0��xk�}��=e�x�>	�
&�vi��u/31��X���D_BU�.���đ��Bl�7ަ"��"���gWN����L[X�����j�KZݷ�j����w�/�%Ed�cl��q�ث0&IP����v�u���3(������S��<�h�)U�ĞX�OmL���l`�/0%h�i�D�c��r�|nE��Q�T�\0���/��yܰEڤZ�8ָ N�U�I�@���l�-�r��-̺��~�r?��������w��:�iE'����u|����Ԋ[���.����T��'��;T32?`哗㘙x)RАriG[Uo=%�l;�L|�n���bR�Q�9�,�5�l2>�����S�9̐�!v�S��t��O��8�r��v�% �dA������\O�@��(�T)���Ig�����𸝜:��N���2T&�Y�-�����$�v�@�En�n6&	�a<�����\|/�sm�s@c)C��ե�(�fp,������㜣�In:r�8���l�,�'S!�B�Ƽ)|�[*aF؂�p˄Uy��ұ;�}�W��6�yn?���b.��;����7]|��?{�͓}F����g�e��R�����e��m�N�kH�"�{��k�6l#/�Q�h��3�tY�=�O{%���/�lU�P�T�bQ�������z��[w������L�藎K�]��ի1ߓ�u�@�g4���@�5Y�6�2�j!Rxib�&L��]!-������~�b��R�
���烋��	��z��O�@���+WRf�f:}��t`�v�����̖�~�l�<�K~%\����r�]�zՊ�ou�rΚb���$i�z�̔.�W7��x��;� ��4��\
A���R+�K�k�8��8�4k$��(����[���kY �mۥ|C%�J�Ϩ�!f�1J�Fe�|\2vޭ0�y<�-�[��3���(眯!$��i��B�R�����`#D�9˔c�q���Q����\�/T�ȅ<��G������0�sw���+��[����D�WRb�wz~҄�T(�:�.�j��C����T�GCkF���URԒ�������i���:<��h<C�<�q��|�׵�gXl����ׁ<P��"�A�,�t�8��R�˄������C~f}FTWɝ��IߛM��O�`�+J>��7|�Jp�v��E�#/���Y�At��|E�)XV���VM���YqHC-��灾>q��f�O�3&"
��������k��j������%��1.����K��߈|d� K0D�$�3nt��qu�'�0�-��:H-h�R��^�f�����Ȁ�R/]_��x��������������rm:�_b���c7�:�z����٢������f0�y�a�w�Z�eψe�����Vx+�Qc���69�w"��:����γ���>mrL0�"�:�'o���+0B�՟J ������o�w	]ͫ�Q���Żཱུ�?l�������0�����{'7�^q��+�`��Wz��r�ZL��w_����ʄT����'��+�	�$����#4����4���)Ƽ��D�ς����x�M�n5r5f�ɧL�>a�;���@��d�\��w��"���)������_�����	�DǇ(��(�{���>���n�2��K����*)m�xS��4����0m�<�B���%G$F��7�m��)��,.��Cѹ����<aҚ�-=��C�\WM�'���KF^�|�Tj���%��D� �����¾�q�)MP�e�<)�η ,Qn�.��"_��l�b2?�|���{�#P}�2q��Z�,g\�"\��xt5��K�����c2]�!�?+֊�F?�8�р֥`"g���r&Ef�+u*��Y��O��d���T,;ߌn�~�<�����Ygkm��T6[Jзvi��8���]n�B�,�`�g�����&�&�*�2�֤p��і��ξ[�)vYf���u?S�l�bإ�*.�Wn[��Q�o��		��+��>Y�E��0ys����5K���~t߸�{O��^�)�9k->z���|��'	��_�]3����
Gy6�=�H��t���`�'�A�#K�b�pM#c$J���a���`�kk4>!�8L�Y�>�łb�LHl����4Ť�5�W���E�R�������:����Z�#�䧫.�{�i��(-���X�M�K]Z��Gj�Os "ю�`f�_�uF�V��w��Dư�|<�T �UaW9����h>����!6UB3h������y@(!BA�4W������-�I�\j�<`C]6fc��_���D�|ř��b��o6�m8�D��Zp�`�\ðI5�(k�+��E��G�/�V���' �MA�#�jcE(��������'��ǡ�=��ל�P*.\P�E�.��&�ȏA2�D���e��O(�9����zu��nES�� ޞ�u%��]s(�o�qVɎ���9[S��О)�:��(�@���+L0��
�^�~T����\����5ܵ��1@�����3e��b]$bS� �D8y�L/��~[y\��,��M��z~ ��,��[��8�a����@��h�?^������SWJj���;���fi;��k�(�-����~6E����q�U��n�o���C�y
�P,�]��ލ�;�StU�O��1~߿������4<Mf��:�AI�ﳇ/�]���-�0&@���pӹ$����1~e}a)ѿ!��������{�>(wb�z􎊎)7aR������ �[�����{�z����ol�������i��(!�w�!�D����⊋�P� �n�Ca�M����%��֋�-���򳛚j��/S/�_;��1�X�ZJ~�rh�0�Xl]���mQ�4D��WZ�v�j��@-�eys�^��9���~�Kz��B�ގ��\�O[�(TC��UZ�|;�6�Y�ߟfx�]v-�|����fa�W*�[�j�V�v��[3��$�~��_��N$�}ْj�V���?N�҅�W��H�H�
Mdw5n�D�55�L��r���BZ� G�&������Px�Ybs�ig���<��]��t�#d ������m��߸��s��+�l�Űe����v=���ǬX�>9�����U)6���[�T/�2�	#��^�w�щ3���0k��R�ֿg�֑�wBK>��o�!\X�}(R�:��R[Q]/�D���.<
�|G��sj��E{+�ꆏU���ŧ�k	�Ir�\%wS��-N�oF,�ˢT����l1�h���؂��Yt�n?�w	��ypp�=������mW�� ����kFIx���V�w� ��fF�:�s�r�_bG��Wr!��19ߞ��/�\��	��2�-�{ɡ�ڕ�v*\6�B|���M�hI5���x��b|E���w�~�i	2j�L�-_���􉢻�j����^F�Jq�� )�H<:o`�U�͸���KDv��.5�p��s�P#P�ҹv�k�#�zԷ��ψ+�3r�C6�8�w��VzH�m���B�3%�ѯz�zm��ȋ�"`f*`&�α:�/���;#q�0d(�AB��	m}�3t�C����& C4�0w�s��5w������`���8{N���>��P7����B��(`�=��ϰ�������n�4'^�g8G���Oo�d^w�i�1B�<ӟ'w:�+���H�R`&pfVL�_���:��ݼ�x�©x��<����I{A��d	�g��=�D��q�����a���V�.�4����`���e�kgXQ[�ԏ������{k��%�پ��e�~VDy�Ś�JL<���md=Q+G�A�o��w�#u�c�5��8�?�hm�ގ�S�imر����a�j	�[܀�yЄ��N9����ݜokNh�uw�����c�^K�O��1f�d����w���;,�9�驨N�ʧ2�1d��,C��xbtT��B��G�4�~wH0D�Z�i��gL���e�b���|���P�y݉�Z)��O�g��V�B#�zwCؽ�T�[�u�X���cmOα��:1	#�F�{��=�{?���G�(S���n��l��Al�1s�F|�J�q/����2�lN�|t�jk1��3)'����d�*'�͗�!'���G��Lcl
�14o�>���w�X.���~�'Lś+��A��l�S�&%)4Q\Bf��ڽ��X�̠SH�6AZ~0�K����njzث*�jk|�!%OZ�/���&�٨�6v��A�aX
�a��=;,�����2V�A��-���/�0e{�;���骞|�!P&}	�d���%s�n�nUf�WHhLgy�"��2m_
SijHA���}��n���S*Z7�'JLGcR�/��a��n�ؖh���~����w¤��Ʉ���n�J��\ԁ��Se��w,$OHS����mߔ$^>D��3oj��V�A|>�8� �����=�)W���t�N�'o�`AL�;릷��xeV�zE���b�x�8���|=�"��Ѐ�}ʱ�`e@�>�amX�5�WK�1�ȯ�P)?�u���I|���~������p��i7��[��oJ4�$Y�i+� d�V�� �G��g0p{��U�����ѶM?��.�U�[ǲ���ķV˱so��f]�ԗ�bE�iy�
�S�r��EP��V���у��ޥ/T�st"n�7��Bh!߫o�������{	nP�w��wPt<*c�A�>�?t�mQA��)#��yZ|x�nI	�q��T̟U�޳�����������ʙ��ZfeB�����J��c��[�n����cg�v~6�N��(�5�f�5k��{�JO�Y�wZ"=���m�c���_!F�%O�2�W�s$�GX����S���p�ӳ��-K&�F�O�����A$'S�5kj,��|�!ơ��O	�{_ˬ̀�h�v�i�l 5-��������AxX��|oF�ӯͣcL�fu��!*s��oj��1`���D�=˹�r-/�Q���OC^�4A�KI�����8;�
zX�mB���g��
����)5�"���fz���(�"z� �27���qiӠ1��7E�*¸�Qu'��O�K�E{4�׍	�6AO�̨�?Y���<<v#iOp��tZ� ?k[t?@'�޿��y�#) _ѱ�β�P�T�YV����nw�:A:��#LomT�����VA]ƽ-���s�R���g,_����DNo��ڴ�j��z"@"�I�?qqL��!A�ƧP��횎�0�|��w9f��q�Ne�e�D���Ɏ�����:��bop`�{�uF*�6����]ڻB�6�.��w���Ie�w����a'H���*'3gM�!�}��ܚi�fAB��S���C&��g�{����˹gVG�Tz���Ҟ�C��X]��ǖ?'� th3�$\ԆK�`�O�
!-�GX�`.�$�����YIm[W����ri;�=lc��ULnGi;y�ޓS+NCϜ��9PO�]�hXy��ֈ"�̦XF���Z���!������g�@���2ҟs�y�xQN7�� ���d�Ul���p����z��5��`�_r�؎����=��Ϩ9p���\2z~�;Ĳ���p=��+!���}���H�~�:�A�O�Ɇ��#��fީ�/y��/�|"���S���g��b�-�� #��tTN5` u�k�u�d��6e��󅫽��@��2�a�Ԋ� �aYzОv�_h�izvg�m/�Z.r��A3�c��p�vŞ�d8��G�dnaB%��4�F�W���0}i7��$z�-/wz�^��-����lQ4a���D���!���G�S*rҒ�pl����m�g��EP\[��z��ӷ-����T3-�־��yͮ@�E�w�b��
K��e(�^�"��.����h�S�݀���"6(���,!����E�6'Fo�;���8A��$��5}@xWk��&�$�*�y���yd�)R�WE�)^@��_�F�驨���ĔG�[�mK�r�6n���=jߦK3���$���Fg��^~�)J�$����%2A���0�A��R&��҆F���@�?U�ʩV�"_XZؿ����伺��)���UN�$� G�Y+� ��[V ����|���F 1f]z���0�Jk��Ffg�KR�,�vo��'�f����c�����$8�[��Պ~<�k�p��O?�=�a�SgF3���s�~�Q��p3�6.lF���BT�A�;a7T����I�1Ul"�vr^	@�ɑy$@5{����|�C3�
v�y�n<}�~w����b�6(r��W��KM�m�h��u6fJL�z���W�`\�8KD��E0�T�3�C����'�K]����A���h^=���lZ�0���P�a��8�
tq@W�Uub�Or#�S�nN�����25%�CǺ�5.�>�7�Ͳ"�y|�����l���?��VB���9�AS�KG���6/�d�h���B�4�?I��b����%V���t���0f��Y�2�3��!�0�1�A����h��H���"B@(�#B��=C��p�U�v�ŀD��Q�?t>qEi<ẕ�}Yq��v�������{��':ԱN�����\]:U������5�8V���r&�6�&��d�P�@�^Mc�CZ���J��q��
Ͷ��gJ'7���u���GY̓/�ҕ�	U�!z�W.U��L�^7�M�3�O�ޝ��۹E�_��`�qi��'�ת).�9w̮R�g�JQ�坰�btZ��o�(&5s�_����Dr�>�sȥ�����u�Ѝ+iLݽ��ֹYV�=g��BvLv���\�,�"Y�7�Q_$;a���?,������@|��	Y���0��4�+�qЩ�h�sLF��e"��}���j�W"��[w��]>ܭ|5����ں�� �0�R����v��]�������*�CLsW�*�֐`Ԃ��c�ŷ��S*�ѽeJ֜�1�3(�Jg��yU�6O_��t�l�G��0N���.+�!.7��xbL����;�ym�;�	���.��翯rЉۊ�}tө��F�,���*o�7�/ika�gn�L-������A����^���3��M��
�q���q����O-��8D� Kﱧ��Q:�%�a�(	�e�����\h�2u0t���8|�2��&&W�{F��Z��pu�rpb���֩�g	�����q�~�e`�86�g��-k֜@��>C�ӫ�s��*	/��2x(���пޢ`�XJ��\U#T�j-"r��t�$ͱ��D���φ�K�U��g�ӄ�>�ߑd�p`їf��%�F)H>�Jt0��B,5���|[��5��Y�M2Vu(D�ɜ�*�Ҍʺ%9-"�l���e6�����'��n]_��P3���*P����Յ�8s�6\���W�Q�t�s���K�����i0	vd�nC��4g��f�Dl��&3���&��JLN�uQ�{,��?�L���'S�D�޶����U��'�v�Ѕ!U�O�5���Vn.$BM�u�6�j�IȄG݈��Y������R
u��j�ql����n�-T1�풊��0�S�r�3���W��>��\��D�?B�&䙵N�m�����Cx%U��wb+���g��6�7HmZD,
S��<c��,�1!��HH���6�&H"F���Bٵ<�L�v�E�1;3�C{�.:B*�/n�Z�B�5�x�K�-�J���x�Tc@ Ӟ碽���je�X��}e��<��8^1�Hw����k��OB��J �3!��>e��.(��V�w�{����Co�����J[Vv#Q��,cFus:���B�f�:�'5'�����h}�t䀪�	�����	<��R|�©pX�'l�$���<�&_��v�l���F=���#�x�JǹJ3�lڃ)�̔q�>x.��gws�WoЭ��u�}pa~�m���f�a�I��?�L����.��F�׷ߑvd�89��S�l���Q]��}�lF�1���A���m���K�I^��ALX�b�Rܘ�4F�nM���h����+�����uR@�f���K�
�6�ַsT�	�R��K�m��r�D������#/���{����c_D �p���2-��*�q���kw҅�_K��6���B�����g��
�AI�>(
����E�>��nș&L�w
/.��27ks���}�C��^��Fo�V������
��6�7������f��f�zS.��{��tǕi��,�!��6�����﬒��G�n
5&�������z���*T׫���<�\d�ڪ�B_S���S��	�����i��ߐw��y�f�)_���.�x#nt�5��2Wr��G�9���gǋ�Ct��*;��.v�M�0���"�ꟊ��,+fG�J�4C���2�SmI^n6�$�P�e��C]BfM�mkμ����&B���)^��,DH���~ � p>b��Uώ�^�74� \��בzE�x�E^DO����%�,�����������Ğ�K�麀�@����� Ti5g�'i.V���zeK6��T���B I!>7k$She�� ��-s���ƈ��4&�E3�\��Y8����F$= �J�S���F��/��Z��^z�G��w�#�;�3F��F�X�m%�K��Z��c�Z�P��b��#6k�bS̝E��T��)2����F�z��k��
*D�69.���uĭ�������|d�.?�Ќ0��.�K��!���-�&Y;�O]�c��y��5CИ�K�Jy�h�>*�\�qr;\���9I���y&@r�ߌ̛7K~�O�G��SZ�PQ��\4W��q�����k+\�}C\Qpl�٨ �x����p0Pd@[5:�^(!xq��A���(Iɜ���I,N�HF�v?b-�2��Y�,��N������D���_��,>��I`:��O4��qE�w��9B����/tr��2D�d}4�a�-��5�i{R�ԇ����
U����c���T�h)L��S���F��.���6#@3G�ܥiM�$�%�6�����"o�o�e���G��g�P���c;k��_0��q`��M�n��#��TBR4�l��j��J-�'y���HU�X8�yXt�l�m�!*��D�s���|�WXFb;��k&'k���g��D�w�bzb�{p*�)�������&>�ִB��j�����@ �@1���{F�:/-�DE��.��J�\������"���P��:�F���^%be��;p�w���U��Y�ؾ�i�Pۥ�u����q���Z����,��oY��<N���o�a�R�����`�h��/S�2���l\���	Xӌ�l�jg�[n7",�ЩU����l�M³/#�#�Xs���w��b $G�� lߚ�gvq�o��u��Gy��^l���^UF�� �%g��'�ؓzp"���/�8�J�z�����I2����N�nXe��9��'��JD�Ys��`��k|��y嚄���+�s��3��+�ʣj�3��XD�~�K8�8�s��i��&]�A�?vI{��c��Ru��&*|2(���U�7�q�����k�q�RZhɊ�YW{:�-���eİ��w�c�-T�\�/��X����Ou1�hb�x^5�I%�����ÐCղ�7h�-\��1����d�]��T.�^:��:Q `�'b� f��ͅ�����gX� ��(g]V��,7�O��B�儌�F�?k�|�����5e+��PFG���׃o�j�k<e�0�yo�͟na��	R�jE��;�FJ���ֹK�4{�֮x�W�������5Tb��9�l�OXh�3�(OGp�T����+B�_P	�-qU�~�*� \'�+@�$�l��8�6�D�~�z�7B�����6cge�Mؖ�=���K�1�� �(d�$�lbƋG��@��W�_�ɪ��<�t��D$��><�((W��=����B�\f�x���.�	�!@��P8MN�c c)w�8�+]���|����鲷�s9��^p��� ��*I_%�dc؂<����s�R�&��FE���1�]�:�K��AW�)�lT�]́B@~�k��uN}�0���Yh! �& g���);��>������V�� 3'��؃�pV����07�:�d& I�>(ܻ����ل�V�6b���0���tB����O8��(>J��3s�k�?���˨z|�������z��<��+���<����~�e	�6�1 =�^z/<N8�O���ّ�:\�z���G>��
N��,��^����6�T����l�����j#(T��g���0�#,�gm��{Fu��>��͡"��QO^��x;��ɠ�c3�n$w�0�2-�x{^&��{�/����O�:�Ѵ�)O�GvU���hl�b([Uur�4�bb��M0i��C�-�t�@5A
�Md9��p�ؾ&�uE�_8��� J�`�i<��/\����z+��ԓѐ�p�'5b5�F�F��g��7�	_���մy �6�|"ϭ�2 �Q��u�*o̟�>Ӫ|�[
�(�L��CY8��٤�q�NT�a�U
M	�p���@Z����>�-�oG�V��J�o7w�����+7��[��}�(sUc��	����>z�t#��r敟��N~oNCr�Ϟ�I��z���3$�]k$ohJ�gG�ԙ�#���	�*��0*�F ��?�c��+b�d�5��<��9�	�nQHyV�!�hGT'<L��tڕ����F7�G�P�Dǽ2�F96��XQȀ��������-�߶{�c���H�g��G�~�<m�F?yz��N�&vg�^�uRzɶ�I��f�[�ww��b]�_%@96`��ߌ�n���r)¢O���$֬�}��T���Y�V�O��T�i-�1���,�jw�pу-�Zk� r\66/[D�����U�2o��8ȟF�i��i��4%`e��>O�[���6s�O�R��!?��h]���Za;ݻt�$��P�s��K�;�Q�7aR<��֣_�YV޲m4�;�؇�>��|}/&�r�<��Hj,�.����f\�+��H5^���Y��F/D���Ұr��3��)��CMu�k�J+(�W�@̸KqmL�D%�y?��-�e���mF��2ߨF��'(���ݍY��p��;Oód�f���Q0�Z���5��Ita
-~�G�'De'�rz$�ڀ������	Wa㭯_�y���*��a�a(Q��ލ��/bV�lT	���Jf䠪�
��\Р��"���-E�e�Ձ�I�E8���^�ϕ:����>hӱ��v���(wǚ�@�as_�ts��̇;�^����5SO2��b�3U�D�/r�(�R	�+��T��&ޮn�RGq�$���gC��xo]\D�����+���w>��W��ǍG���r��5��B�.>k��H��B��:��ٞ@�[ �`��<#X��LA��V9��k�=D�D#��!�"B�=��/�A��\}�B;��>{����S����ت��,�?�pT0O�İx�^U	s�����es��ɢ��NTgR�����ƽ>��Mh�Ļ�"R�|�f����f�w�y�{~m}��1���D,������5γ��]�~�ئ�X��g0g��3}R�k+��M
�+
�o��Ra��c�~ �6&
yf���r��߬V��ss��,�R���3T�hL���;�~S���2I��a�a�=��D,���n�$��;�����)ZV@������'�Ey���'�Z����������ّ�)Qf�
!�30�O�mO3� |���3��Ǳ�N�0U4���X���7j���<I/
9��E�����R: -zlo���7ö6��ћr�#@A�0M_���ބ�����;	�(s��啔P�ٓ+����t�r����rU-t��˽�K	mj��F�1e
��u�X�0�^#e/AȊ�1��K
_rԅx�@w�#�"o�6��q���ov�y$�q���GEG�N{y�͏��۟u���_c�4\[f<��_���L�n���D����[������4qv��/�̥.�a�/�H�l���ƌS?F�Hi_�p-pЖ=H��lb�5}{��� 7�G�+H�jQ�=�3A��n�ڥ�D��;5�:�μ0�C��*ʭ���_zܸ[`ix�¡�Bej�,�MpY�z۰3����A���§������5-h�xJ���$�/~���!�m��R�%�P���C�&>�����~q����T�Rhz�Hh��M+?������|E����ΏH�����#�2` (�ĳ�#		�e�ĠVsç�� ���8�W���h_�J �+Q���bi������[�nv��\QA���m@9m�ɍza�o�
URaf��si�f�
��ւ���Awj�LB�ď`�l P�5ס�Y�*�ڴc��9)�p��fiu�����B��[
�%A�lDp�=MFMU7���Y��Īz�V����Y�%,��[1l�s��$|5�VŁkf�|�a�
�FޤC�b��h��z�ĳ|�+�Fe�6�On��p�����
��\����A�,�D�����:�2����}ւnO�/H�Ve�G�%��{��!tO���Z�J���,4Hd�w��O��a'ȈH��ܒM�/�h�F#M}"ۓ�V��k3�1>��ၜ�f����,����y�g��5��8��NL�~|.��E���3�$0��\��	�S�niq�qq���w뻷��xP�tDxk"�vA�U"Q��d餡�L������A�T�)۰�rF��0_�eg�����lx���-�!���p~ϱ$�T�3:zr���i��t;��y��3�N�KeJ��� 	����Q �*���MLC%��	�F'�������&�j���ٻ(0���W�����4f���,���S����0�ܚ�y�38�O�٪y�G��\��:���I�jr�ؘAM]>�� w��A����V���hr�KN�`� �����$���M�Ig�\+��
����L��i�|�(υ�;u��� >��?��2z���t\ r@�=3b�<�m��䰽C�4}#���Z�LZ�&t*���(�g�a"�Z����}�]���2��w� ο��rrl�q�όv�EN���YF�g�����]N*nK�/�B����3��2������E���yf�W-%~
x���*��ʄ�ϙ=t���5��~b����׀?D�*K���@l�,��@��-Sb>�mbz�Ƀ���ᎅ���ſ(	̯
�9ڕ�O�"[l*��.��z
u�&=g��a��V<�:YN� UR?��U*GE�g�������I#Wi@�[w�P�*�DF�׎+�K��*��	��\'�=�c����׾���3Lث��T�Ә��ƞ8����?Y�Z*.�!w~ ��\�t��9zm\����e�������	�y�3�^�Զ�9�=�ASC�Ze|��L��6�͝������f�R�!OH����)G�y64���0GR.������fĜ��_��^��OA��E��Ca��y�O2��$t�!_�5�'$`�ET ��"�;2��؂�Y�Ƅ�@7[v���0v1�֔(5�UZߔ��w�T�`�ϐ+T��{�=����%٩�:YV)x_��<�X�����T��ֽ�-2}�I���s&`���-$͠��bGJ�a۱hi�K�2�^>��V��V���D��x4�-8
��
�[l�,v ��!< �#��S�L1����(��k��/�jBQ��lO�<S�K��ѭQ�O��J��/%�9�0�����'߻�F*��!ڿ�apX�6�I�+�8��#�����9�N�~-���_�M�?ÿ�+�!�۶a<���sϴn� 4>����e3�[T�g}�E��cMWkF%�]ϻX���[D��	��i'��u)��'�p.�K�sP����]�\p$���N>v����/S��Y�p/B��v>����%�j�� g��$��.������q�M���LV���.�������TS�`��<:^��xr��8��օ�.'5`�l�p��<`�� ڀ��ͽ�/'>F���gNS��N;}@ e����0>�X�~Sp8�W:��|?J��w]N��4�Y+���m�٦��u����ѱ����f���:ZȮ���#A6&�� ��Y�3v`1�����9�+�XupZ˿�]4��El~��I0�^oq$M��\_v�ƫ"�+To��(������h�}�޶}]�5��\�V��_�	Ç��8_8�i���|�߽=	Z��� �,��"�w��'�q�X�а86ޮ@�I���f7=̭�f���m��1��~&�G�g�t�#v�;ufRH������o�
��
;�{x�$&f#=p���k�� �C�T�%�׌��X��7�	١&jm�̰Kjx`UhB��4o$ɘ,�-�XJD�'hz�.���I��\�QZ��x���'���E��w;��D$�A$ #0�Ei�q5�Xtnׄ=n;Bd����A�Vئ��v"���k��b|���ϖ� -�7���?K�S���B���wA���zr%�v�����G��G.��D��+1�~� ��u*ԡ��
��k(��eX�a�����:�� sE���^��G�l]��h<J:�2BFw�1d:OfD|Ln�1�b�Ǘ�c΂JG���T[����ĸl-G���!�L�CX́�1�y)���I��:]�m����m��as���,)E��P��;����
�����?��A^��E��#�b�\��"�Yk��Z�T7~�󀍯�e�9R��h�>�����0��D/�b9�n�Ch���U7>�7ʎ�
��A���έ_����*��ӞԺ~���'D����H�}��(�m��ل]׹f�
�$S.c/���s�y�1�}AHpP)��_L����A�S(�W� X	�i��ˢӽ�:�詪�D%UyRa������<��U��D�]������6��V�{�������M�B`��	�K��M���g�G2-���Ė�&8�N6V}ۑ�s3N��x��,���l[�Y�ނ7����{%v������Y.J?�%Ks�R��Bl�Jz�8}�}�������ɩ8�x]��q�5 g�T ���פli�~�`��f��`�R`o�:���cW�'KhG�1��r��:���mؼ��gL��x�N��ɜ���5���"��q�/.��T⬂�ʤ�c���N(e�SM�F}l��Y���_A�n��]����QX��<��浺Xc�ݻ|K���M(�1c=ʦ9
,��K�8
u^�V#�\'o�C���ĺ'����=���8�D쬿ZV#S�QK!�t��CK��bzW���u'�� ��-�����\7S��ı�L��:������s��GжB�|�8�ڰlB�"y���s" �)<��<�1lJ����~�i�_&5^jМ ���&*>_�<^b�<?w��7�sU���`03��5�\�Ӽ����5��0�呲����|F滮=�� ��S�#�H��r��y����Z�XV���"�0��=Cw�;�חR �(To�X{�Q��=�%�~��h����&R�xF�k�����1��	;��$���0�B��Rg��D�h�ڦ�{�~��s�V, |�۔�CQ�x�wk�W\�Xk�vF{xō�هX��83.�e����<?�-r
��=t����u���;������'ӻ̍�EGy���Um�m�d(nd��Q�f�j��C��@�y�%r�2�نOe�4Ň��*S���z�V�uiİKX�'R[�{��{�@v����D��03�-��P4���f�PG=g�{�:>v:S Qu�6!�Э�4;V����}�n�ͪ��>&n� �~��䢖��G�:.�%GE��x)6��÷�c���z(W�O����j��� q$ܗx�՘n�[~�BJ�*ņ�w����bO�^>�02�DA�Y��I�<]����>!�=HQj�u3 ����A����z:�S#�}���/�7��3|�bL��uxa+�,6�Y�ì��P]�?K4��؄_}i�'C�U͠A�h�Nm.�v���Zj�@X��лWf�}����ڼ-%X��b�b�*�2�灂Bd�K� �Oŗ>R|��T8A%b,�e�Q�I^վ�-bɄ��
P����L>4u��5wOh���mA���ښ;����ӾJEA���T�$���$�%=w{�	,d�>�fZ ������%�k�Z(��\ն8�|��88���b�]��8�"=�NƋ_�^���0g��QY���"	��ө�}�ᆾ9�u|ь�,���w�,[�fԄ��\?��І�����/���gw"���rwErnzt��;T�CV�����[�ak�g�d�O�����[�.Bσa��@l�Td��ӻ���Q'�J�(}�ܗ��W=�=��;��� ���;�2-��Kўk��A�BL	 ���3��H�0����ڲ兗N�!�������Rd.?��BJ 6-qur&#�;~:�Z�`�gUEw9�0��[-J2z��:�3���$aA!��*�ڝU�z�Y��,ɇg��GF0
����bUu4o�Db7�s���l�O'��du�����B�m?V��bٛ�)NWW��'�o 3�BZ�lu<��;�a!� "��C���u'[�\�8c��h��&&5J�蔭�e�*�{�,o�
6�F%�@����9y�
�>�0�T�<Ďߠ���ɿ��gN������]1G!�f���4Ć�e�^4j|�6s�x��Ր�Nտ�
ʰI��KX�5���2�I�`����z@u�M�9Յ-@�����.<����4�P�Es��>����zb�`��6;����1Np��ʏ� Αp��H����F�a�y��������1�E	�" 1�ޕڞ�7���U$�-����(C�c.��ъ����u�{�u��|檣|������4�|�S�O�|��S�IB4�!$_��!aA�z�l���K+yQK-��,�w/I��Y�k;O���)�*�l(��0��Jt�`!؟��JZ)�C��z�2Om�WRw>�q��8�<W�&���o�0����+�p�j?���{����BK!e���X���S�mBy���r�����V��u�i�ͅovf���q��]j�)A"�S]�����H5��J�P�pЂ����=C#���w!�Z��B���b-�i�����y�m[��WUOe�s�UUr͔H�yJ�"%~�*�����s`��#{�.��k �E5<��{�?�����9ݺ<��B���8t�$kv6���(�uE(I
y���J�6�`�^b�SFaRk�qϧ����=uVZ�p��ʻ��O+O�D���>F�/n��Df�G����'��'�������-���]���.�@�KW�:)y�W��{L����<eu֠}���~����^4R� V�y�k��t��9�vyh��ϐ��8h�0��@�6+����ï]&K��lhM-O��+ᤫ<cs��pӸ���)�5���G{����E�U�	��}<�Ow;I�m�\.�ۙR$�Rv��V�*���.���G������{m�(�R3g�p}l�����;ʀS<�b�ƀ�l)�y������g-!�;ڔ�r�j%�1��/�.蠈� l�C��>0���j���=��G�IW�mY�ԞZ'Nn7��c�9� �kN������SG��~�~|�ijQ�\8TA�S�T�icl3�h3��]����*>�����Xir����&�T��"�;�,e �����Df��[��9Ki��,�ȫ�*K�[�8�b
�����$�Tn��ZL�@Z��HϜ��T�u�>ݐ<[h��x��zg�L\U��2_�\@��u����bPUw;�^͂��q���l	�5F�V[-��~Ua�⠯�V0Y,R�E����V�df|8wvG�,�>�w�=#2�T�]���B��	D�J��a��xq���;�#�-kHb��*K��)�r�Ɗ�	M���Ȗ����F����0�˴T������	�0�Q����!�ȜJ#�f.}N�}]+Ϊk��E�M#2uKG!���p�葕�|���(1: ���tR�jl��{j!�c��Gx��w��8�����d�o�f$�ֲj�փ���%�A����
��~����+��'�%�RϑHH����A��k�K��I�{��0'������#���!����8Ɲ�W�į[�i���p%>l��?�ڔ>6X��L�T�^ꦥe�F8�#w�۰����k*�]dѩ������+��z�P���F)HU\��	@"zL_�>�:���,��S�*r8g�ɸD	��Oc���~��&w��.u�u�%t�9� @���Q�V\ �D���he���8���+�	��g�mWf-�E��
�t5�u$�U�3��(l,��Js9�	�EQ���.\�%s_�"P�4���+g`��	��1!��ަ!�s�������톽�Y��I�1(=��A�Ԇ�tM��D�zי*~����@�	p�
T��洪z_w>Z��0b�T#�b.3��.#��n��Ǎ��T�(0��ę�o�3�6b5����Uz ��l�Q$�g�g�'��[?yJH��8
(��C*|c7C5̷$���mIgg=gث�(s����5��]�&_vh�D����k	�^�����%͉YJ�Tb*�W|��8���G5���B��"�Q[��vNG��E1���KAKJڹOh����$�9@ZeݘALx�9Ï�6W�sI�m�Z����K�Z����gP/�y24�:(J�R��.R���_ѥ�W{|���/�6�}�\�'6&O��.{�G���=���\_��l'���1X�˹��u�������A�1��%7�I��-�>jv�p)0��֡��
��|w:PW���DԹ����Ӻ8�U"�v$���^ ����a~�a�Hd���[A��BH�&zл�!gvA�z.o�,O�eOH�)���<��+j��ڄ�k���]���X�H����?[:7�"��1=��vF&�c����~S�|[8.��p׎���>�H�YkC
�s�^Y�qck{G"�����=�uLh_�+2Z^�ЄG�n@��P�P�X'��}�'L������ls��4�|؍vHb
�r�e�wq�q��#�ɂۢ75у�19��2֚�W�8���-A�\��fk���0����=f��u�е�B��GNѝ����-���Xu���m�!P�
�v���*⏒�:�������S����w���m��XJ�5u܃�4���en7���̵h}��R�=�"���MM����~k3���� X��0`wn��GSɯA�R5��/�E�oS��E�>I��Ctk�FB��uQ'\N�� ��e��ݲ��E�SGk���q��1a�E�$����*_괍�%{Fhd>��!F��9�g�[0>�������11n-c4È9i�F��wVsfF5�u�ߢ�\��ٺ��00e�tڬ�΀W$��gw����$r9AL��^���I�i��V������{b����W3Gx��![`^��hFP�fR@��7�E���A4oS�ѧ��:c���G��ͬr�na��R�z*�A��'i��֤	U���Sc�]�%`�@ɋ�9ݔ�D�9��Q;[m�E��Ls����g�g�=��J�R��;����F�jsk���G��[��B�G�lˈON���]iǾ����P��ܕe��"C]��VјxM��R2.�#��6�E3�{�,ڮ|6��4][b��B��S��5C�mܓ��v4"z�?��uٮ���ӀD*�㎡��{ F����c/��?��4��i'��[(��:"GJ-�~�<����ť��@Nq�T��80�6�K��������/)W��x�pZR��8pl��<��"��	@S[ R��e_&�z�J��	OY�ܕ�g�Ľ�딙���'�By�������3E�I���%��L8O�����6����A��%v)p�Lү�!�y(���nqRЭB>��7w�bXk��ps]{�uo��"���	��~��W�S�q����_����J�CLR�\P�97�U�4��kØH(�������΋��~y�M\.&��6�e��w.jlp_��GE�|$v�Zd��i��y	�����Q��B*A{��]���-��g&}7�����c���!�{��?/{#�L�wRhN$O �e�%̧h<Y�mߵ��8�{��+��)la��V�k�	|�i��.��u_���Au+�'.�4#��w���J��ϗ~�O�x��4k�Ρ��;��eo�Ӻ;�<y:p��s>]�2�9�)��<��^����h�/�+t'��>Q�@"��V�����"k_��E�q\��A�Qt�4��	��1�v�\�lk�)4��(>�_F�.�8�L��D�A�����:�1!wIU���]�ݜ���k���-g�\�MGk��U|�ƃ 3`S�s��3�"f��3c����m�0ԙ]���u	�_]�Fr�Aæ�^���:�E^ ��=ȩ�\y��։J����a�m����^Ψ��ɲ�x��ٿA��'۸�-�^3;n�E�,[_j���̑�0w�]Bk咉��Wڤ��I�)���Ҷ���by�0�A��e�(F�ZL�G�������U��k�S�W��D��zr�۝��|?�����ֶN�}��a��r���[��rǱ&X�ǻ�BfZN/�6YM�Kʯ��8�1+�qG��&���	7�:驶���S���������:�������ό��O�n��G�fj��<K����*����7�1��Y��E�9���-�l�[؍�;��eF�p��#�vD���b/C��E�lp- cR�ve#�C�Z_RK�e�0��`�k���X���i�k=�0�����7.� ��[kh�ج�㊊f곘6��m��W�Q���cFB��;h�EOUK�bpkܪ��V�ߔ���� ���7�����=>���E]��3<y�~��"1 h79"����%ݳ��0	;g�����;��0�ngA���;��a��Ǟ[1�j ��.*<||�e��r�C�F�n^t'�10����[~��v�)Μ�ƝC�^�͆g7�7�0*P3�lG �e����(g�O'7T���j��E=G�h����. ����L
��ѡ#��W�H��<?������a'L�j�d�v����EK�|�DQ�ؑΛ$.Pb���fX5&�7m�{r�� 	��2~D��B<s�����̗�8�������N�qY�s��l �1����7�Z�G1���[���7��b�vч~X~�J����)4)�YJnw]�yJ�WU��`<+C3�Օ2KZYl,�j��CzjK���J'se��Nnh�}�H� ��t;@�G~D1���OG䝏`�B�HWϮ����uBe_���u �G�Ѡd�!4z7�v���޶��E�=�@���#��2�h��y](k� ��$֌�^zy�O}�Y�k�B���Sv�0���M��u�2y᲋��A�CY��iL	kbg�=�@u"���a��֞SuQf�H�l��M����#�1�����>��lc[�G*�f��Go|~P�b%���;��8��8A6�h���α��'$ �_},Jу�
'tb�Ѭ�z})Î�VU���C��ؽ����d��A�Q0�h��c�A��E�\L�7GG@j �zT�0��G��F�,Q��('��d�z�YuGҏ�����ԫ� �Uss���%FE7���s�P�U]�:�L��t�5���!����nc��I>0��rB��A�ñ�ϐ���%6�����fx���͸��*�6�-:��Y���'}�7�]]=�qmd�s��θR�-1dK�����jh�ia3^>�p)��n��Ɣ(��XΒ�����=��<���E���4AD��]�ci���t�����0�
����;�@��_l7�jW�y��[fw�� ���JX���bݿȝ��h,�A���_��v��Y���D�S4ċ�Z��}�@�/wz���;��~nBb�zȸg�]�C�$27����ݳ*�\��oU��玕WQ{8b�^lV�2"��L'��R�Ea��݉/:}�ĩJ���@��ɇ�2L�}GN��[�9�Ղ�,��JWhϰ��8/x�X�����}䵞�}ٓ�T¨dC�p�CnOc�-������Es����7[R�R��8W��".� �� �R�!�@����M~ ��X� e��f�`�s}B9��i/Y��Ä�	^��o�E�'/:e��ySwYW�dE�d�k����r�㊝FM\*����-��w������eQz���?(�FL"��?J}�V�-/,p|�QW�5c�!߷��	Wn?�����Li�M@~$�����M�h\��_0C�0q�	�I�`��b`�
Y�%8���4�f���|p2�y��O�4PS��cɨ	^R�0b^oVhWќ k#���]�#�^��>i_Y\����BaU�F#}�����d�"��9�������I�h���o��ba�u��I��^Ë��!�k1o�0T<����1����9�c�3i�P;�Pp/�.3gV��p� �CN�?�M� �K�Q�E��3�j�ߊs>�e�I�����HA�p�>���!�%o�U�`�v�ϷN��~�1\��KD%&�@֘�81�D�r$ͭ$@��[
S��,W&�q��&�c`3` �����M�nj��!uw�% �?;Y�˕�f>Vl��H#?�����«�=���^��L9j�zh�Np�f�iOYQP�=��B@yҶ���#�������"u���˖��p�:� �����:�Z<#-x���ANQN<�]��4����y6<�7�,�+�˪�]ٷ]�ѥ�Ru��'�(d����z�W�`�ͱ�?���F�\k�:+c�$8@�j���k�����0��d)�74�X`�Wk� �b��o�!p���QE���o¿������6 �}�x�;�S+mLK���vބ#��wU:��$��6vpi-�d�y,c5]��[�Ǿyٓ�8�����-;q]<�/ˑ���DU�8���$���'m�Z\C�E�+z!b:	���T�'ꃍ�]|K����s~Î�H՗}4����-H��Vcv��{�W`)ĕY]��%9�q����<*�˰�vx�(C��K���R���Aa��ç*|�U��sW�r���4M�Ԙ��P��.�0�1��z�=��d��Ƅ�����K.��w��g�E�E4�l	`fk��T�)К��9�=���)�2���Y�q��FF��,�k?$,��Z�R�F�;g��T�3V�X�h5�#����W�W��J��4ZZp�r�)U�Ah�4)�xŖ@��Qş�vPA7D���r��>�0cv�!�r�j������Ozg@"��w7]��G�v|���M�OB̈F^T� �y.�S�8��� ��|�Oy��"���8~4z�����`�PiI���f�З��[�C��a&񑷨�Ӂ]��5{h�Mb��f�"�[�;L�8�r�T�lEg����AU�%��%ude:�ȑa�"ҝ�5I��G����a���ư@��$�}���G�t"|���促F� Cu��wxq�C8l��.��c#`G�]F���M��hfˀ'X`¹5t��
���YӾ�+���sЈф������e	�� p5��?.�-�2�#�I5l4�'Y�ϨV4:� 
��\9g%;N��-�`� ӈ�sh1l`/�SE߂�/����;��+�!5p;�BS����v�2��~�a�c.1��Fj�{J�F�-��>w���y���Z��ڸ��t�u<"�k���#��Ce��B�1~[����OjW��9�m<@���Ž^Y�N�S�T�|j�Nd�.�0'�(��ë��Z�y6�8���W�i�΋���^�SJb/�]�d^H���w�M@�r��z�NAvO=ΞV��@$*n�?����J	�0ߘ��=h~�(XKFC�4�0�_v���i�����7�D�6��%�?���oPsc�:��R��4Hpz�TE!7�&$]j��d��L`8FˀD m���W����u=�zN���]�a���c(Lh���X��~�w�,��:0�*�13��[��K�Z��xK�*���	�V���A�(�N���j��A%ƴ�1n���,Bs%��;1�Otqf_A($�`s�R��bx�׏F};*|'
h���N(N��p}UiԶ6��W$|�-N�Ͻ�K�tꄚf��~�*>�RBa�a⬸Q���{�ʾ��,Ϸ���a��	�!c�"Np�}�vU/�a�T/և\���jz������w��m1��ؔ��M�H
��T���������*X>2�F�\뙋�O�<
M�2/��K	&@ݻ�?����c�q%�}ȿ%�G��S2�ƐH�oh!�9ˏk��	���G����zQ$~�0���+v���������A�ۓ͓u��{nl�"�]�o�o����2��Qaq�l�A�������gU�Rhl�p������
XM��M�LP��6�od�2�m_�'�͇z�?��1�9�,��]� ����7 n8�mP���;"_��� ,��֩���7�&]ڻB�[�jA����?(^��b�s�$AZh��5-(�B9��g��C|�y�ʑ�s|<�֕���X8pQR�F�0�����MB� m+��}\p�PäD�y�	mW�!�E�ޔ�U����֔���|���x&E�8h7)��T�`�я�e$ܫ�nG7m+\2�R����γ��8�:(���_�ƃ�ڶ��}�SC0����@۾��6����p������(�Kr����%Ĝ���$�TҺ��YJx��7����_�JM	ΟF��P�V,�¦�2?�e�	�ޓ���*60��&�0�	L/I�B��8����|&޴��/���$��N���`Gl/�<H���g�3��
w��?wW��F��%{$�I=��|?�>�g���%OQl���Q7CE�wq�|0?�}͇(g(m�>�"��5�}����?�
�ю�'��q��]�����������e�b���� �B2�U�s�X�v�	Fo�{an�҇��:��r�w�H���2� �އㅱF���������T�m�jE0��7#������j}5�%�q�{�xN��~v��R�Ub'�m��妏���~�65n.��J��'�|���?���9Y��Y�7a��c���G"�p�C%�Ҏ���Оq~:�<e9�R�nr�p���<�� 1U��>������S�	�r���+ W�tD1s��pַ�<�S~+J߉\�,�����Ajn��RPގd�p�R.3}(�|ٯ.���^�> �bm��7�o�uV�|[P�]�
?XY��V�ܕ _��c�-g<�ѝ�_]����^�}:؝!��0[�O2`7�cEQY�u�j� [7#AaP�M/v��u���p�=.s�ҁ�/����$3�b��p�h�]^/�Zi&qKpE酮�p�j��p�2��X
=�)J&�9���CS���7-Wqt��u�ކea��	^x���d��Vc�f�OEMy-�G�ܠ/9~�ݤ�[!��bX����k�O�3��ٷ~�Ec�F�MS�[s��g����Ps�Fm0��@�Qu���*觗v霨V�+�4��^,����~�Z�W�|t�Г3^�uЕ�tu؂%,���Z�?��Ԏ{��*@��P��M��g`�-'���3��cnafc*���ܦwܷ����<��LP�MAK����u��0 ]:I��IT#�n��}O�}cҬ	�ֳ�"�̿o���\��R�'��v���T�ېA�a�+C b���f���+��&F"��b�Ȑ�Z3�R�}^it����ls�C� 淺���bZ�#�m8��;G}�R��l����=k���k�%kOߥ�
-��Ϸ���"-�z�z����+�Pt���R=ҫP���)�q�}an�{���x���HWh=��lq�ε���j�g�n�ع~�;��R�D�@4s�`@D��*����/�Xգ�FU'G�L��ۺ
~�����՞V�c�JMqi����C�5r��Mۻڛu��,���Si����	a�^��a��(0������{�����^X�	C-v�q쾚" $��QA�	Թ��5:z���-~E�4`xE*��`hn�-VDb4��˻O-))�Hq7"���ޜa�+�4�6x��+�G+�7i�!��t��sp��%r��_�j�M!�g�S���f���w�)�����q�*�J�������h��AFb	���`gz_�)����>,J�n*}���N\��g#���;�荤�(,���{:@G�8���t���rL�yp��V�^���� t��� &��X������6}f�SxW)؀p��!Ə��W>��7'z�RÐ�K �����������2��5�yCdε�Ig���v�ʘQ�c����@aQS���C�F��j_�9�,f��Uh��Z�l�č]��.��(P TV����?�����>|a*��I��?n�� {U�A�n��c�P-u8��*�lu���(q�\#��iDc��������TVƵY'�{�n�!��)�s^��7�M��g�/~֘J � �QQ���6���hug%͖E��kQi���&��$����Щy?<8�+>���QZ 8�Վ��m���^?VS,F4�6�Q$Y�#�J@k�IY���'����w���T��dC�]�j	�V:@�� ΍r�߲����v��4����Ɵ�׃�r~A
�&��f$N58��vB��?EՕ^�pCG�2�ˊ7��;�Wq�t�_�!�������ϊn�+�������2�*����Di������<v�D�V5�?�d��o|X��D9����#�0���R��J�~��ǆ�M�|`հ��M@�n�*'�1��|O�u<��V���5R���D��2X�#KQ��-(ӹ|��e]/�*���_MZ�x��	ȼ_Z�sl�F����;��9I�������R%w(~+�Zf��g�j�(x��V�L��g��1��SWLo�l]7zvmr�De����xD/�MgF�8�����u�T9���[��9�a3�f�_��(�κQ��!��f��NI�O�!�p7܋Ԯ:�!��f�ֶ|	$�>����0��{c�_G$gNwQ�K���\!��45���h�P�w��9r�G����>F�BI9�*��� q��������%�7�-8��:Ǧ���'�X�&�I�W�dY�~��*~�P�̪��l���U�u�0�2}� �Mc���k��/z�1#3���:����^�u.To�/0���"�f{��>�RfX������q����˝�M��EMmDc��6�<5�w����ｊ��>��d�S���X&1�?�Ke��?�N�;�bx ���L@�(qR\���KOa	��6�+7�Ȉ�D;v83�G{��3WȻ��N�	�4L	A��"��'�)3�wv
��gGQ��Q��b"hZ�M?MF�XJ����1�U#dpt}����L�M����w�d���TD���x��"��-�_�B���� 
�_��1��;���ɾ��~�Y�S�޻�1&�"r<��_~��bЂa��������羥 W% �H��d���ފYI�
]��ek��M��op���꟏#]X��Zq�U
�$Jk�nS�����m{~���m��8)���R�'5	���PZЇ)�,{#��$���k[��>��
�:�Xxu��߰\K�(�������f�j��R3w�����O����C2��.��`�g�o����n!��e�8��1�9=ι�}w����݂���?���@9Iq��n���z.����,0���1�'|��shm>!yp�g�v�@Ӑ$��r�b}Aq����3ѰN�C슦 K���(��4�4B`�G1a_� LÚ)	To,��1o�b�P�DĿ�o�T�	Q����,-dlD��{�|��$����c��*o�_�ٖ(#�ə�{;8S���ޅA#2L���.P��p������_Q�E�:�ۃ�8]C���7�!'2�eڄ[�zr������A5�?q;����Bj�ٌX0$���\�:�:C=��'gg��sE�Y����o�bD�71\���h�(m�L���I�G-IєSu?������0�Tx�tKI�h��eX�v�Jt��݇���`z��������Ky����ҥ�G�,9LE*�ܷkw����-ϱr�)t@�YJ�O�8����o����:UI�V��NE��9�D�S{3� �]X�e���X�4��;�����N?�l7_���E�@h]�~���Uz+p�M+�%�;J��A��qpt�݊º8�LhUڭ�-Ub��3�2�߳�]�h_K2�ޮ��/j*��(6՜��z�j�Y�:�S�gE
C�����R��~�?<���7��p�:/�H���Z4P��Z��XڂW誝��R���;��<���*<�h�A�ֆ�0�fT�{��8ꗑ�Ui���s]㦟�^#p5��He崱8�GXU�`��}����-�����o�)��Η t|�mW,D^���w*�j~��0I񻣶��=�����$�쐏�E�mk
�����������/��5��/W���i��9���V���=y/���iX�Y~�ˋ|�ʶ�5*�� �0�g�eտ�aCԚ{8�5��|9`B>"W��/�]�D���k�\7���(�ɹȴV�:�����>��ܬ�p��l ����%�		W�A�~�1a����0&�W�<bz��\M<z��A�9/wK��������P�"���9.��;��5�S5k1�1�x�y!Ĥ�#6��Z�"o�_�(��Zef�-��mu�䷕uv@}e�qH��)��W&�S�{���Kl�v]��Z��#0x�����W�8�IN����	�)��δ��]5'�)�e��z4]/��a������*v��� A���zN��}#Gӌ�>f�T�)�or��!��g�j�C�B� �8�_v���G�?�MW:[֘2�����3%n�]��j",$bC ��H.�c�o��2h�'CC��V�E�#�V)�z����z���:�t���w
�Ƈl�jm��Q�bk-��J"���cf�� ��H3I&ؿ&���FT'|���F��ե���`䏀Pusش�&f��brKO��%e6�vkԡǱ�ke^+F����Mڸ9��
���[�og�&	ؚS����C>s{d��O,B�i�n���\Ί�*q���<����M��g����-/�8+[�=HO(��.��C�6*�P�K���z�ݣ�D�@��)CJR����\�Ȣ{�ߪ�dF&8��6,��8��=�D���EL�w�4~�Q���I@7�s���-H��e�a@]E�P��=gC_�kuF<�7�ԝÆ��q7?����C6���ڙ���&"�g� K.�8s	gP�礐=��pH�j~05IT{+��6�s쒛w1-��
�@]�P\��� V!Sߎ���s�`�(��%�;W���|��~�|Fm�`>ɇlO�.� s���W�`J7�$fz񨁨�e��R14����R{_�~� ����Rd�0�b��C4�2�@����?BEi�	�w��XR�9�XD]�4 ����	v�_0^K{��K�-s*	�Z��%��ܛ`3�O��Il�-P��%Һ�(�W�\�J����d<ѧ��6ѫ~��e���0Wb��<���}	�/�jd��y��|�1�Mt
Lv�h`�����=�@|�[�H�)��]cd�Z+�ƪ��hdd��e�§T�|�����.!`��sHv��}��1�"���ǻyC��������:/�L�''��V1 �_@�i���N���Rq�Pj��L��B�ō�(�7��u��2�l�`���r����l�.�V��*�cܫ� ��l�z�����5��J��}���ێ^D����R%��*O!��2��щ�k
����|�lm���Y���-�y��2��y�e��)�N]��R#H�x��ߝ���R�C瞶sHnV6��֠� Zyd\����ꬎ�iT�e�i7�U�H�w���������f�@hs��-����zݍ�3�^f�B���,����n�4W�V�s�@�G��dЮ+���WFZ�s�@*��\����	S�q��o=
�^N��W��u ���4@X�΢	P����e��J�K�rz�8!5�J�t���o��O7�]o}yM�E� ���}R��ì�;F�$�]̫6�O�1�2��e�|J�l��qZ}Df��P�"xEG�u�Y�9�D۶���#qm���k��]~L3�� ��;�ĭs��c��s
Ъ���H:�K9�{�"a.I
}ţd!Bl��5?��C1�I�����3�ju7��#hk������_)r+3+��W\�Kw��h�S�z�)AL�����#�ҹ�>��?/�8C�;��0ǊRT&�_����ٙ����?��M����Y���%$ɣZA*�*�ţ[��dY���)�N^6cZ;�Gn��r��҇�_F���^��!�v�{��!TA;l,���Z�!yN�{���Em�n��������6M�9U��#a�;f��S��:��|:n��/]R��v��o*G������g�����@y4sD�N��jkz�]ժ���8Z-B����~�Y^v���ըG�DIg[[�'�I"�	"�&��Cw�}0sZ�&��@��lza���G3�
4r��X�
"��a�-�P����4�n1׋�ӣ[�®�%���**XLE�>td�QJ}��d~T��ȬP5&Z�~����/�ʊ���ђ��6:��	ʁ�����V��ɒ6����\3T#���I�F8�~߉�w�:)q���8���"�V�"k�C�M���枦�Y�μ�����'��2�$xR�F�o�,�)f�(�K׶Z=@l��v��
6���Q��1/�B�L`)�����B��r:;v�/סC2�㙃W�I�h��Q0�:$��'-$n��f�M���K�%�bl/�2����A�^��`��6����8h�!��l��՝�bU�5����*��yԾ�"h]wn�%P4P�܋��fg��0��g� 0:jNT��6�1I�Ѳ�>�Z�{A�|F072�8B:;�j.&;�Gk�6�������S�-�c���y��բkO��De�+������f�m�� 7md���n$��b�.d<t��S�Wډ@��OЫN+��o�6����4�G�r���Z]��*?�e&CC\ 'f=�o�Y:Q����C0��S��6�-�L���)�����὇BW����-o��Y�:?��W��,s�U����Ѝ��e�ã2�f�Q.-!B4��Imy�z�9<��c�H`��*��-Yz�d�>�"Ig��¨�It-�®����h>]��3�M%?�[MƒcS�j��QWz��$y�c��<���.n5,L�pJ���+�eD|��%a+͈�M�c2O��
&DA|�S2%�QSF/�pTs>���<����6L�V�5+�^L��h�VOh
3����H�$̤���C� �$H���B��j	�A����i�e��!�g<�ڥ��%.%��<�8Z��S�����+%!a2�����z4.Q�3���K0:{�Y9�j�E���a��}x�v��/?7���N���c���С�F�j�v9�U����@{��ޘ��ݷ�+���YE|��۶��k�8����-U-PS;��[��NV&#���_*/��(�R~��Q ���1����~ �d	,˷{W≡)V;���ݜ�E$����5�Cx�ɏ�A�ё�7��	8����!�'���.yv5|5�`<����H6��x�&�S+�2�$�of�XI{�u=R��i�p�ru�IY� x����6@��vӇ8��X"���Ȫ��������V�82�d��	�M�"?1�C�m�@� j��B��?F�@��ӚD4Z"�-t'�\��M�I�[��iP�����4�ñ��sk�% [`��"`+�mO��qW�Y�R���P���m���ɇ�{1���\7[���Q� o��K������S(\+�]#��:-W}"�pD ��/P�*����C.Y�R�*��p���w�pK4��p�iN\��y�9��^�o��(��)y���p"�nRd>EJh�[��h�&/m��N��`$�E�W�N�Wj
ǳ
��"�}|���1�~fԣb?����}��7�y�Y[��aN4l�������-� ��kU��;d��4ڬ��L$�]>��'�|�Y�?g���c���F���/o�9p:���_s3E����� � ��W.�^�<.��ۨ����ԫ���\��ewx=�
Ua Ѽ�'�+?s��C_o��Jyrv�۱�WGSf�B�Iz���ݰ�5~��^c�����3�E�CFEݐ�3ϗG]�|9�?V��eoR���R���X��@k�`\���L����ڳ�дTL�3��N��	��6�Y�ѧT���a�<�U�\�l��N�j �NPn�<NO��hl}�l٪
��M�&_\�9R��=S}������IS�M$o��!�p맶W)���7ļ��۠�h��6v�%���єe�����w7�u�vdF�U� �.�Kي�h�B4��0)q?|2��̩D��N�]�_��X9(ʨT�q�tC4����Y��g��\M��G��| [ￖ�,��N�0 ��)��/��h*�'�1Hr[�B-T}ȸ���Ο0[0ђ�2�"	�I��ɁV�q!$ڏ9&�p�k-�.�J�kzoT2[}�R= I���4&��p<<�5C�i�Vr�ān�%#V!o:�!`@��6��s8�ǹ%\���G��e?��wA��������#�Q5c@]䅀�tRF�L[O0�7�	�:W�JhiHZ1���y�0�&cۊa�Z�1l7�p��Z-=Q�2Z��gaB�*0]�L�,c5��*���E��.�3��)PB�7�=��2�KAu7跿W*6�!q�	�3n�U��������l�^8�@��lݳY+w0�CF�|�>&����fQ�%��Kx5������T��t�oxa{�O2G�`��ULh�Z��z�N��� ��*��jR��P�Nu�o2$�iet��K0��t4������E�E.�������L<���J*�o���g%���3 ø�!aJ�T���/�4`2�F�h6c����3謒�/%��R�q���}��E��.P������`P�IKrf�c'�\�wM�.F�1�ʶ6Dt@��
�.UL�WX~�^����T1�O��ɸ~\���eP,�@]�p����+]�>�(�Ʀ�9����O��4�K�T�)U�"d��GC}+��W���>��N�cS��Z�ܶ����w�f *��bN'��3R!`�Dx��2ܠ���K���a������\�Г	���ܤ��>���[����/_�'��oF[��ƺ���>�`�hyQB..��}�=]���]��AI�!#� ���>/'��<�Y�W��lb2봄_#BЯ^��sf˧^(�:԰	 mC�1D[B���FcKFZ$����U�K��ā�{��`Ƭ��w販�z�]{���3)*4���H $lj��[���ܠ��~� ����Z�h��9�%��X��3�ý�otS�!"�ێ���O�>�K�������f�U!�)���G4��m�N�SGx"�K&{�:G����Š�����q\s��|!r.e/����Ý���ο:�%.y��,�B����U��~"���I*3�I�K$ƿ�;���1l�����to��#	�7a�U
]����5�.q��P��t5ԯ����q��.�ev �>$)Z�}~Zț�p�Т�w%���т���G��
À×���nb8�4��9�E��g�h�L��FH ^�b7�bI�Z��W1��C���R��ƴԿ�]TE#���_f����ۂ]�%(�*$�3����:�86���#��:]y�?ԨQW#�_��y��?����5e�7A�`T���4�
f~�������|L\��W�Z�j�Ⱦ��a��� '۪�/��yzf�ut��zD@`�QD}�����'�f'r�f��I��h�xP�J�л���Q�O�B.|�>�λ�7h�E-d�	2mq�;O7�ڍ�o�L�����^:�Fю�Ak��Id{;�=�������<��
�c����Z3q5�T�EUB�RJ��tI�/GP�\��9�tD5̓�dX�J{��c���+���G��1�	d ���H����Vb���Ia4�ṽ�-�&N�=��6�U�Ԉ�ޓzK�[�4p(�c�C�*E6!������8V��&+<�m�j�-�|P�	׌D�P۟.E��!	<9��">OU�ڙ$���`X�o��4Qp\p=vl�yihJh������j�C���d��G�%z8%��F<;c��{�t��~�!E���)tWL\׭��D��n�wV��聈���j�)Ͽ�E�Cܬ�
[c��l��ڨ� �X_&K����$��(��#� o�n߅9���n�16@���#)�Y�@��}�!�����}T�W����$ǓZ�B@��IȰ"�R�<�B��jI��-c���{\b�s�|+TP0R�P@��vO����"�G�	;�գ�����̿�e�Xh�M���S�����m�.��dkO��)笆v8��f/qD�KىslSO�ҏ�ie,C:#�+�a�J{Y��W ��/�;}t^���c%��ӐQ���9�1NK-4|
�BBa�͵b�sB�B���vk
���'�b�е;,b��\��9�Y��͂���y��̤�`��/��F��k;G-�Tw�o4�%NE��_hzL�y)�O,���J&Vޠ�`)��@F4]e'��
���qɵ)\(�K#��Y�74�y&C�PMw�w��օԑ!����Hb�ՉnBߔ���lb� � ��.j���K��Q�Z+LR�A!�L`�d㞷�-B���_�A坂a�p�����&t�:4����8�>��n�������l J�����%���Hh�=��=
p��Ĺ����n��|x��~;Z>�@4�L�䊜Y��D�8|���6�g�y�,�VZx����<�>���q�(�c��$4.Y�>;���/�$�j�{��b���ɷY2�hq��)��I��|{�������Ei�9�"#���5)�`��.�j��EOFR�R4�+�W�,gt(,	�-��dR�c��Ԛ,#��A�eAw6�+��0ۃ�����` 8�*����6�����+���!l'./A�SzϹU���e�vA����މ-�ĆT�0����a��d9r\>(��v��WN�Z����ͱr�o�V|���(l'�͟p���U3��gv��@�A!�\`�l9�E���f�>�;�%�lb� �}�s��-���G�o��Т-w|iJ�a&��G�{
�?|�(�D\��1}����h��u��9��+�Ki霣�xjY��M��"��O�v�K"�yD�# ~�&�8p1a�T	�n�Xj�U΀ļ$,0�8,6�@}G�d��ap2��/�5��e���|r*��=�o=�U�;6�>s��)�'��8u��X2�&	 ��|؈�$���gC��F���4�;�.#�����>�*y\;��<�q��`��fYѡ=Z��An��%7R,N��5k"�-r��f�n74�v`qs;ﯼ\�����o]��!3�/�,aCa���?.�P"����O��J&6�Ƀ*u3����i[��@��n�4��'ڀ]�#��#�1�b���O�0n,dW\����*z���3Hr��֡�3�T��H���!dlw��<�P�!Yr�iY�q7�J�ќ�d��N!��	������Sb�3��rO�����)��8�-}�5�(
I���>�sb��__�r6�&�6P��qj�2�w��9��C�5�Y!�첛�;�Tb?�ë-KK$�`}ixv���?V�b� ��0d=��5��BA͂b��*^�b�`�	~A�y0)w��tli���.ߦi�CUg�IF��l�ǔ�/���7�h��6e�j�"I��o�y�`��h�5
rp���De苗	�ʼ]~�+��wL.�S;ݭ����hT8 L�����~��/��%�o��=�} ���H ���>�n)��_�h�JMa���WkLU]�(2_W�\X�PA�t����H���	��n���"��a�kq�`B���8�8���B	-��s�-�
���ңk�I:�ź�蘥N�j��y�\z���i��@�&2j�=l����މ�e�������%�7i90ܑ�g�]Y����X2q!�ӕQ��Ȥ��MTj�ƳN��\.Q�f(.��;�-�����N���c"�' ���u��?�A	M�����^��'N?���ԏ��Q��ڿ�MA?	Y��.�ͱ���1�<.N}���ж��S���#�nq���o_�S|6�Ej>�Ɓ�-�vIE���~g���$���2f�x�'��
.ް�w�� �#1
ΐ|����8�0����bZ|U�M5�oa��K���[N0=�z2���4�>����y=3�+�����f=��ewN:�]��A7�������;E��	]1L�7Ǳ2;M�w�a��	K�b�Ճ�P�u��Eb1���
_F)g��KPjU�z�3~@E�e��cf�F:�;��RC����WZˈ�Q�P��д���>l[���srg�M��e*-3 j��_�x%{	�e����湀�͑Q���́/�{�̜F��sD���nȡ, �ƪ"���E�!5����=,�M���3/$?EG\��+�;�q�C�b:����0��Nc�DM��*���	�h~�u�u!	2�6�`��߬�H�?W_����97�賆Dg��B���t{e�T�	$< ӷ�|�o��6�g�.����
�zAj7A��c4"���2K�^ɲF��=��+�'E�@��	�G��O�s�nQ�$3����MDM�ղ#����2�� �M�]����*1�X��p����ѱU�$�j�pK Gq�),Ĳ���������]̶��C�;�귺n�M ����<T8\��骋���u�����G�3S�:��j�9��V������!D�8zp�ɳ��M��4Xϴ3/E����)�^�sX��\*�L��P�87 �!λ�Ayo�:�yZx$������v/楮ݍ�j��Gb¥��HA��	�-�k�I���f�:�ɬ�գ!ٟ��21�ђ�"	�``C��ç<j�:H;�x��a�ؼ�Ln]]�Fƹ��8d�?��Վ1��(�~v�=0�;�O~m�D��Kx�6�sL�07�#w���!tJW�\.���
��_���O��8N)��| ��Oa"YZ���Q��լf���l*��0��}D����\��ןLj�vr�II�L�B�c	�cIu�0z���>@=�N"�\Pr� }n�c�f/��HÓ�}~�c66N�t~K�iS�.uy�� V`ʎ�������_�_���L��x�v�8B�Q�Ju�E�� l�v�$o�D@ei�8���~�w�I����Op�����$�)_f\�ڃ VQ2n9�1CN;
^��#�1vU�ĺ�v�jv�m�-i/��)�n[��5��x��Bor��D2���eU�˾��bE�a�Y�2�c]��nA�ɫK�>��<tTi Ĳh�%��P�n�C,���L 0�y7�ϭU��zK�G�Z�U�"I�ou��%���ۤ������܅�¥���//A�R��w�~`9���5��ѿc����$�0(<ʵA���n��߲z��<�M��_���ԦذU.�����X^w)5T���i��yG�D^�J!����=^��YOxQ Л�:5y;[1DY��J�4y=YV��đ��E�@+A�߄"p�3�G�w=��V���)��(x��r��|<�ߴ�,�6#���d#�K�(�����/z��a�9>��fķ��:`�E��O>�λS}l�Q�5i䋓����Ǎ���1Z�&�uW-䳜B���A�e�]�i�u���>V�j�&�&�ɗ\�2�E�F�.3/~)BP��3j����r�2�hP�K�fi �D�m
�>�wL?e8㹫���چQg<�b�$���rK������is��'z�0Z�Y��=��!(4*��3;nCMWC'��B<,`mP)0e�DB�T_Cٞ����_�tB��7�̶<c�5kB�u�.�[g�/Z_�p�����o��%�wB�ɂBdd|����IDS�
�`�NZ�:����jKzy���NX��J�~mr�pC���qz�7wf�*�a��>����%N�o6�������5�O��^�<O���Y��r�ڗ8������T��cA���mS�F���t�����G�r��qr�ئ���> �a��Ӏ�!�6��$�l�?��3��?Is[n_2�A�3E5J��R�Ui�z`+��r��} ����̀��~�c�?��	k�8�^3v���s�
�����M��� ꅼ뱗��Wkdֱ'K1
9��l��5�P�����:3��e�pW��}��JJ/�-`~�����|`��_�����J�������� �_�}� ���Ū�����Ĳ�`��U��
��<��~0��	������i!S �� 6b��K���R��IjZ�^'I�u�B��1��� ��kM'�!�̧����]y��[ ���ێ��K���(/2C����g����"n�,���_��ͷD�`
��y�Yp[9��d�2(>s�w�0�pǼc8We���yv�a���<lm�]��*8���n_��B�!'�nF���|I?��1m4�
�V��`P��|�la�^���I��=;��k!ː�Q8*��=��l��t"��-9k�X�"~&1j��S\A�t�OF���=C&�.5�?������J��Bs�W4�܈]-�"$�M��o3�����<�ceorx��2%O�����u�	����!�|o�2�Ҭ}�d���+2���h1Y���u�#�i��t�	�P/	mX�:.�ŲZ8D���֨�n��}?jb����!�W���cu<!e^~��R8���9u�/[�}k�S�^?K#�i
�C0 /�.���A�´�wz`�v/>c�@����:��1|�U����Kv���-�9ǚ�M~�e�4�.� ��i�l<���&7�+���Զ��)z"`f��}�t3�r�Ed�άJ���� ���2Bo8�����H��aA��j2�x�@�-#�|�ധq�e�sh1�ظGC�|�d9�Zp��a &�G�x�É��,����]�0-�����r� ��i�e��$A��5�Jn��xɺɑ��ޫ°�ܼ[
� ��'�Z�|I�F(�0��c��"����8���M`(�FH=4s|Ca�_�1�2^����l]��;j]T�G��x��=YIi�[]Q���3�r�/,!9��Z�ID��'ʫΥUW���>6�u�J�_"�آ����Jj^�!]Ei��Y���X*���m��Z��k�P^�񁔇������4��|=F�[9��x�H�ur�����e��	E�\�~4A�v��]/����|7�w��R05�Xb�a��b�Y��0�Pȯ�|R�[Ii���sə��EM��%�2�(��y�QA��*&�./��������bbj 7co� ��Ggr�)��μK���YAAO��������dMru�&�Ӫ�O�De
:P�1:6�l�U�����U�s@�iג����Ni���m�N��	���P��Q�kh�JJ�`[���>nM?�&3X�p�d��K����[l<�k�*�Z�	��l������CY��s�7�BL���1`6�L�ܗ���Dek�&�@Z,��7e�t' �C2��X�g9䥻�4�܉�7�4=�l�MH��O1eZ"\�Z�Y$�+��pl�q3��T?�+�oIw����k� 3S�:���R@��ǈi[�NY��s�Sq�λ��� ꇧ���渫����	>���Ѓ���{ �BYޒ|I�m�L�x��n}5����W�/�3'9�������c�EV�ED$)��9Pn�̑,0;_�X���-6�a�p9����s
emP�Z�e���o���NJ���H��
t�b��{O�7s �DD%���W��X�B�gm�����JUTX��|=Ih}:W6��?��`wW���e���d��������;�E���t�w�M?;>�+gU`�b�ׂ��ڼ2�f�/dz8�h�|���O���kׇV,�qT��/4��D�7�؟���)����q�ȐB����)- ����/^�'���n�-���(� F�~?L�$Ъ��*rV����jD���.˗i�����ZE�����)�r+��z�f�,<C'3�*�^;��}�c8��9�":����c�t�򶆹^6|A��e�{���~$�ځ!�b�xl�*�d@�QG�et�RY�;~5=�z yO�\`(�)��$�?��Vp8��G࢒Cݺ�w�i���zu@HF��ǩ�h��c���'L���Ν�Bs�����yo@dD��+_b��<�O~����i�њ�{h��%�HjT��?��x��<����X�!ݏ�-�����z��2v�?��GU���	��4NL�֚G��Dt�4ָ�� <:f o����u�g2��"��8T�0���C_������T9pw���5=�'չ^VR���PU4{�{��t��� .�a�Ẃ�LI/����[�DCH�'��s�|�*CF�:���}�7�k��1���z��u/��Xh�8�)����mp��!��v8� vw�y�a��4f�,ϟ �{�܎�@;�ld�΁C��Qr�#�6���neC;��s�mly�[����)�-g[������j���\�1� R63��!�ё�[��.�_�L�{�}��oP��`"�9�_�K��^id��h"фLF���8ٖ3cԛ��3_�*���W)ƃr��:?�Y;-�]5�w1�;oj�l�x���(��z�nrtN���\��b����oU\���9Y�R	�ٍ�S'To}��P��JT3����Pa�N�7�h��܋'���ә)�דm6�XR-@ߣ�KJ̶U@͒��Ӻ���B9ݳ`΄ѡw� ��5�?Z·�Fj����-]�}G2�+B�ވ�vy*��y_aIy �[Y���B�4&����ʉ����42�o���0$ T
�.�q~e���J�en��C�FiZܫU��9��ꂁc��pқ>�pZ�oϴ �c�}R���Iu������ �;�i�;��K��0����?�Yiû�@a��AJ�O	��Pa!��)�����%S�F��x�G	4��|����,+ÿ6o�zOVn<��1Q��qH�z9�h˙��"{���22��
6e_"Y�&�n���
_�LV�2-1?Z=?W�D�:p�o^?����a\+Y��&O��=��ɄI�A�+��/<�A���Gv��f^�q��8�< w�?[(כ��cV�'4�����x��C�XsR��وl 1��uryUǵrV�2�8�҅�*�#��lQ�J�>�,Q3w�Nt<Ķ˘�I�������CU����y
���y�B!(��]?�mӲ�:&��Ҽ��8�O�����p�6�gr�u]J2����յ�@�Q�zR�\Ԇ˨A~�^�^����hX  |LSM�$L,.��K��b�m��Bj4=�"Q�l���#�����2�f�k�����9=2E���BҦ8�+'	.h�
���y����}!`�'�OP&L���6��
�����QL�l�������/uQ���-o���#/�4����@
�7�@�9��X��ԑ������a	-7����������H��5���<�oX���{ڤ��,�����<-�N@a,t�e�y���@�ɜB�%#���F�:�\ӕ�.A�y;��+����ԩ�(��L_lG�6?�|��\%����'�X�������aؿ���Ģ�x�7������ �ǀQ�}(�)��������E[Ҋ��X�
W��8�4Gt��A��K͎z�=eD�����wf��?e���{�9۝)��eabsV_25�u@��Wڈ�6k�y�*��|�R���y�%�*}z��;�.�����G��P��e>*��n�[+�| ��{*�2���{G&O�:5KY��֞��25�+�1#1�[��Z[&Zl�E���q+�������Uo�5�Ґ�`�.�	�8?]M��}�p|�s���0�'t���AS�Ff<6�I��D)�}��t�)*����v��}LIv��B1!_��I�a�ޑ&	~º��: �A�I7����GJ�3����s`aB]X��}+��p�3�%�dW�7H��v,b����ݲ!����ݵ�YF����t,���d�sxz>;	�H������=+�3��-�'QΔn���}�����@_�`�:��`�W�SL֋�\ଆ�x-ǚ+ i<������d잤C4/�����|iv��E�0~`�T��mI����PSƾd�ɷV$�Y��{��^�H��=q���?�u�xw��R�Vf�>��w��e���s?��¥ģra69w������L����4o1�����Z���u���~�̀$wާK�˜�̮/ODot��w���B����\<��E���:�����|��5�����1	�6�K�VXK���?#�ϼ�ѭG�GH�p��J�z!/�?�H��iH`�]����rՂV���磊�cqc3�#��=|���l-*7�-�,Y�^�$x�Q�P&����l�`NaR��0�A�0�ׂ�d<��ܯo�~��XK�3ҕ�FPv}��:�Q�H�W����=�C���C��Ґ~�T�ξl����zH�����E|]-	�f5[K�Ohl��4g�������[��ؕ��W�k����hy�V���di���ݏ�d�%��A���o��}�����?����f<e]F��!k
�>�Ut]��bݺS��{D����³h�*c�&�Z��]��O���D^ޓL4`�	Ad���e?�uV���O0yW��M����1�����W�6��{�Ǆ���M���Sʬ�RCP����xUv�vG+|h�R�x��ja$ � pJ�S�Kh-C����/F�`>�
�N=h@6�W�'���`��>�v��$���&:+0i
�k��V'=����'W1qیZ+��휌��4*�Ԓ^=$��U�������~(s(k�� &�Bxe���I���ּ��[�,�����`�r�|tm�mD���X��iO�Z$‫�`��I1Z��Mip�wS��:wl�.��2��y��o<�c$y��U�&+���n�����B~������W���zO).��{�̼��7u�O�|��kȮ6.�m5'�P���Zq�P��q��Ps��ٙ&�}TM�ٽTj�y&t���n�T�"�m%��$�n�φb�Ejjm��"�vzɀP�����d�`���8�v�h�}j�<�l^5Vؗ�'d3�1JEוkp�ͼ=�γc+�����}���z�/��3�B�h,�8�R@$?tͮP��'m�[��3T���9�n���Ki���}���oN�r���\�����t;;�esm"�r��L��h�GBX�HEjV%r�^2�5��zRJ	��\��η2�F����3�5/V��)�N^F��6��܍l�Ys	�rV�ƅ�FȂ�*=����x�p�l6DJP�Rw�� �r����M�C������*7�&9���`C�E�>����R[�d/}ƽ�1��z�j���و��� Q�8Uqj$�*,=��8�A��]�(��mDҋ�n:�&4�/�Y�:t7��!�*�}���f����k��&c�s�eg�-Y���	�ܧg��藠��a�{ؙ]��p�0���N�x��vAԬ��;�%�F�C>C�C3�H$Іi�AP;h��:���	m{��� NУ�FY_S4L�W�I�ПR��k"e���6�� I�*��S��k���Ҩ�/��N��D�^��5!��^�+�)�L3��T��$�;@�PE!>0G�
�[�;�yգ�X��Ɖ��)� �&�����<�w_q���xj�@���y["ű얿m��}�H��$�u�����@�E�î {h�����*p���s�E�v,5�c-n�f˼���=ݢ�(KQ�D�~̑�(��7`��p6��iV�Gp/�ro3�ϡDw3������;�'9��5?�WM�T�"��?�������D��{���*�yw�H�����-����T���Ȱ���<�x���lv���� 5�qW��v�'s��&�~�����k}J8^�*�i���R�-�Kf�{�h��n�,5,S�hwNA!�,�G�
.��ɰ �	�a:�X���`?4�0���Ĵ��&��`�<J��S�\�Z�U0e�J�7���j���	�h+ڞ������]��MrY���#�p�����G��?u�?|�47y*�f���=H΍b
g]�C����|�M!���fJ�BD��֩��V�hs����
]b�T"��W$�h�L��R�cc��.z�^h,��q�}���
j��B"��~W�"�&#vPҨ�3�&�x5�l���-���,H|\Aj��#zm>�� �������n���J��oy�2���A�����A~w��WfÃvv����.z���,��r'�kT]�Ҵ��!�c�a��/48��CŠ��]X�2RL���8��ÎZ{���f�_�0�PC`,�4��~�)�h�=u���Go���/��\���e+|f�\� �����>��%GF5%�^��9�k)��ƫ�~%{#��=%K���{���|tc怦x^�z�j*�Ȭ�� �^:�uA��k%_y�A�s��EU�������Z��w���k��h�����%�q5�H�bS��<���X�gm�v;�bN����g2O����+�n�h(��Fh�6�n���q� @,��-d��xЎ���\/d>�ؤ��
�t��p�=�z��U�΋�ܱf�v&L(@e��_l��u����}H?�����8���K�׏>(�O����lID��"�Եy�����r^����u&��5�R�I��	�']�p
�z{��\(�ږ�Ug�W�|���r�WIP���.�}��]�5����G	��og�D����m�W"������R|�V&}s�ly��ePHf*���-�bմ�Az��LE�LRzF�������ޡ��ч&����4�O�uKC�C��J������j?6.}��T)��7� �.��o�~_.IA3gW?g����'�����W��p-� ��1������D:�J�m���O]��;/6Ϲ�\q�����]|e�Յ({�K�H"�%��f� >	P��G]��hb��	]�fM�r+eQ�*|�H��y���>{�ys��?n "UL��x�d��k���\j�g`�YJ��߆�@L�2s��.�{��1]�!�~�Oe@�8�5�kO�W�ӭܩ�&����ү�(��c��r�v��=j�SRcM/�@]��<�y,��!;��=�X��Q'�NT�oRM�M���2��R}k��v�	�i��bk�����.�B0�~BT#S3�0k���k���/��C��۝��U����2��[� E�n�b�Ec���cЄ�P;�9��N?�����-���U%E8����cm�ҟ��D�ק�Nb���.��[UO��V��N�(&�"�g�-PE�GM� �Җ=%p���_�ɰ#���m��0"��>T����q_ǧ�|�gk;��U����Wh�����W% ʢ���mr*=�Iߴ�/������F_�ց�@2�*h&6y���,�O����S�ɑK!Ԗ�Ih`l���j?�T�ox�.�F���-E�1Swe�q�<C��"Bv�&�yQ��x��������T4�����ǅ���=5�0���}Ր��bwC.,�2�Z��j_�'z�w��>qE�����]�rɊT��W�UV��h�����+��ys�K�!�
u��Vojv��'2U�"��&�����K�{���P�9����˕�c���٥`����xy���]+��?��7���ܸ�̳�P�]��Ľ���@�B��$UOH&&8������{�^�kH�b^&O<���$�s@D�G¦���E�)Kq>e� �$d�.XF�$|V�i�\����SOcs/��J��B���ӆ�'�+�p\gYw��/p���&ǫ������*)��{ˈt%��p����j��:���_f�b���V,z������ͭ��.��� �&���H����WG`y��w��%,�.�_'�ua����'�W\��p��J]��DQ,X���n3�b�;�4:c�l�2/���`
�ð��c<�v2���
jq���o�\yX<�ǐn5hγ�W
B�_�NZ��H,0�&�0�����
k@��H��>���뚻�ߚ{a����p��ztB��"ǥ/�}4�d����/9q�� 1��o�ֆ"?��	|㶘�3;;����G�Nj>���\���͌!�p�����c�x�=q=����$����}6(d��3�@`�Up�'�E�V�>���⊡c�	���)��Dt����C���A�׹O{�A���s�Ȩ��r����WMܵY�dTx���b�x�\{�{�n�Gb�rk��7W{�ˍ�,��G͞�a\R�x���M����C����xZ-�WY��_��m��Pkk����`�`�~��������=c�*J���*1�XDT��������?}ʈ�/�wo5?l�	Qf7�e�;iW�t�v��b5� U���U&�f�v��Nx��;ScyOx�o�u�����^M�O'�Uz$���OA&y5��Vŵ�ş6�S�z��=�i�LJ>��>�cRI���qԲ������i�gp0�_kt��L�����H�3���ݿCj������$W���ˌ��ܝ�Ր�����v/�K��\´$3�[C�3�b�]CE(:xʏ�����e��7K�W׸
3�#�9�3K���@B�f)��&}��a҃�PR��}ہ�W+x����YcbgMH}g,��]M{r�EO�ݻ�o����^�C�%�S��qg�0ԕ%Μw� �p���xZ�k��O`��踽�����@p�b�-��|}����G�T�vd���=#�m�G4�MQ{�|�#�В�E"��K�
��4�͇����.l9~�s��Ҏ@i�p^��DIx�L�  .cv?�n�
����眺~�DIzU��(+��4�7��p�q~�#�س�0��T?�i�:,�5��b��pU�S9���񋫬6V�jp���V^&����ɪ-���"����r�Z��D<� �X�Q��-qp*GNN�&"���\��LD���=k���?f��́���Zl/��`�ъ���K_��x]%�,sm;�;�Q0���c�pU7�jqd��:���b�9	�[�����uԥ�����,� �{��f}#@S��` ��(펥�܂ǆ��L]�dl]����7-�#�Y��x���~�Z�o���/�]m,D̽IT��mo9i4Q黂�W�4s����X�=���������-�@����n�����;Aq�%�b��]T%ֆ?J�U,a#`�_�;�0@�.j�$��n� %V��ƪn˛�[#����o�����>���Z7:�	ø&�0��zn)�t�v���rKV##:FݻP&��8W��.�H�~�*)���^�	�eI�pk�̓J� ��f	u ,��.ZL��60	�n]����O8�:��Dd��7�N ��bR�*���x:�Kl�-�I�P�HМ!@��ej�!�G���߲v�M�'��j��[��@BU�u�D���T�+��d1����c.�R�&���us� k)��8E��~�D����r}`a��o�<ԍώխ
M<"�;	qy^�����;C���	���m'��Z3xEl��Y��U<�U1���a3P���.F�-ه�k?���~K����FF�
?�M�BS����V�t2;�R�"�\3������o���g�eTX޼�T��E�2�那�T��%}<n���;���l0�f��!��I\�K��8?���K��0��Ľ�� .0�4��{z�`�K�����J|Z�ü���;�����@##IF46�j����sՠ��"�+��Jp�����#���y[�%Sf��w1��0���G�����O� 8���_
��":���B	�0�4oO�%�p�L`"HG�X�x�ʝ��)+K��.��i]J!���3I`���ڥ9�� �����$�7->x|x����'֊����#�!&�`ݖ�DL��P���ʔڂ��NE���ya���fs�y��^xlV!�@�_�m@_e��):��,!	��
�D@H �ݍi�N�QQ���/�  �9�����(̎
")zN�� *B[�,�����b?�K�$
�wt ��:���w,Ɉ�f� 8�Zta�&�R�q�L91�z4����lh�N�*���m���BR���U��-�m,�Xz���t�dIXf*���|!�.�@-�;�.��<����[�w�~���p����^����_�/\�g�a:E���ND�
�-�]��n�Mb����=��iĖv���g�Hy�35'��4�t��!"3�2���|Y8��fo�le��TXWm�C�#K������+��_�,;n��R��s�s��(�����V��B�R�ņ�������Ԣ����F�'������%�'ag��
���d�E���;5&���
m��d�i��K�8�U�b&��8�w�(ha�]�h�Z�i1t��[�c��dr@�K�
I��� U����4(؃���о|�-�qڛ�/�mG��+
�����t-��f[(���kTP�&�	�6�s�p�Lq�M~���&�H��Ks�Dܼ�/N]4	�m_�޴TTc|�M�� �i�&��f��Ye�VWt�"��/&���|x�S�Ѡ������&���@���o5t~�aꉪ�����n>��i���,850�$�W���5��H",+A�'̈g
3?ct����ي��Ø�%4�,� �u ���J"���]��H�oItd����&�NU]{�N5�@�"����2ðy�������޿#~`�(���}����z���	�޵�	˸�AR��~O������o2��� WF����Z%zU�h߽]2ݜ���5�Lބo�����V�E]~O'^�"3�d�>�7}�y\��bݫ,�a��R�C��:������+4!_�-�X�h�����r���7���vE�Z44I����p��Q�ϯ�vP� ��&�o���m�X���61_쵃�a��r��{?����G%�Q�U<X�*6����SPF� �Z����	�I4k/�C�� b��]Bx4Tx(�q�W�3�!���D�Z�� 2����
�ehb#�wB��' �{�LZ���_���)�K�,>+dI���cCi�C��f�`b�����]���~� [�A��6�T��;�xV軭t���Á�c/��bz��\��tff��*.�;�@��{4�2�G ���J˫F��)4�v��?O������<�>Ԅ�'l�{MQu�b)+���(��vC8[R�ж�Y���)o�� ��B3��pk��U�&��$�-G��L]m�d'�� l�\���h�3[�@��n:eC`iSPf�>�*e���*��W����*�Jk�����&�wk~��1V��=�e��+��ϯ���:PF��w{v�8	����w�2K�~Vzbh���q��Zⴥ��;we(>�
T[4��9����ώ�W�(x)�WUzj�rR�������2���<ߵqӝ��K�K��
Rl�����9������V�ٙ�9B�8k�k�X����r���\��4��E�5=K���c���׾�Mc^�XMZE��ʀ��4�/8jS	1-����j.��X�P�������3o1������(IK�"N�E~�(̂�ݛ�C��gI�����Eq��Qgxy�4�$�*�4��V�T �g�7N���Q����.K&�#��3�#nFFC���L<h�51��|A���d��F�)Z��{	��֝/ǝP�QZO1�$Ғ���3������|����#!2�0���c�����Ƕ�H)��] '\�zɔ���������̉9Eb��}~���XJ����j��&ՁA7��	l\�����}[ے�*�����6+D� ��}�4�b�\�,�pNB2��%��{�
��R윉Ux[Ir(�2�\g�+v{B'.��&Dy�w��7Ҷz�!�X��
�ZF4�ܸ���Y��pj�)��
u�A[��˧h��oZ�2]䤄[��]�0�~a��4�(XHj�}Al�ښ��~�k�b�Vo��Ӆ@�}`�t���Ji�L�" �&(��s|p��8gL������#/����ֱ���������ʾA���Qt�Z�^�A�7H�7vЧ?������f _�r���ӡG����^L]��No�I� Uo��y"1�\�ym�
���g���N�A�Ķ���'V�__�s��Y�d�G��;�S�~��:��Kp? ��ؒ��5IePϡSVA�^e�S�\����o��W��]6¾���Y�d�AzH��J��U�[u@��o�,�@�^���+ڤl�/I�z��Kv��f�ZD#���8�y~�[�W�-4�9���sUv�����[ik��w^��v$�my�؜�>�Ō�n}$��jBr?����)S��2��w�����Lu,�3��0�8��R͞�u���A���b5J$-t�[{B_?��'p=����ly��8�Ś�$��C�&���t����2�iIlR�:ũˈ$�É|�Je3�OF�H��b���UP?�=�^^򧗴;dV�<�B�.|d�3&�J3�[�х�;�4��~��/�Y8�H��E3>*��?�`�.Ծ� 
>ץ���d�
[xĉ/D,Ce�#�B�l�&���?�<��#;k��}0o �\��H���v$A�����-���c÷N�^����Nu[x�[Q�ُQE�b�ి�@��nB+���~x��ˏ �|� �;�RXz}�N�� ����q�bBDp�2v�(O�9�}� 7�i+��^ɋez�4[w��+@���J��	Q?t�u`moH�o�L+���5+������>r�l��0�3CX_���quq�>��������oe"`��q���w�$�V�|�����W��>&8+5H�L�Pt�,�)Mģ箛]��#1���Q�L�!�#ȵ��=Qu�6	�d��
^�w�� �?1#��^u�S*���?ɕÖ� �N�"|Y�5Qdǃ�� LfXE�zU��Է�;ϛ�/R쫻)�g�\���b�P$^}�RK���
�i��G���`l (>����EHE�>`;3���ʿ�A��3�4��#�zf ���IE��ˎY5HoEuO��P�7�
+�����6%�\pI���s���5�? ����|�a���Q�����,UvY�j�cO�������Ӽ����� '3e��I�{U��ۈ"O6��D+�$d���8*yɍ<3o��U�:�p���J.� �'����&�)A�W]�|�[�eg҅���e�>�%��\��ŃrWL$W�����*��.5,�P�,���9q
���a�`��f��%�$�&?�b���!Q�z�Fcq:~�2��b�.�Ι���|�f��!���Iv���r��e�ùj��?9���mB��6+￢�;|�a�z��Q�s��=A��C���)���|�+�+N�M SRc�!	X)9u�ӽ�a��ӭb�塺�Za�-M���#
9w�q[��i�Z�ǉ�f���5٨�J�O�Y��o�o��A�S�%aX汗{B�0!x��!R�EIf$���j''��#��0|���"`p�* �����V3��B �%]h(TIKwT��*)�]�Ȳ)=���sz!�Sıj]p�1ȗ)�Z/�S��]�%K�������-t�����:�p"{O*�7��/�r��\h�՗��ӥv)���F���z�TP/78\���f�A����9��4��߅PXC8�����hz�~먕刾��`}Ko�bX���:g�hI�&_���
��
ݾ��=��7�.�,�`�7�)��|��[V$����("n�ޮܩk]��Bw��!�ɮ]d0ķ� �dk��$Od+q8W��Ǻ��'��0ݸH� �'1q=�g�s��VZ4��2*
�t��7�:�R�M��M�"ӊ�7��]bj�ƀ�/'�<����/�UJ�����-<	�gXB]	��(�B3M��pP@�J�AJ?bp����:_G��*}�R�6��H�R��9I̯TT*Xhe��N���'{�=$����0y����OU���eU+��3OM&�)Ω���C�������P�'��6	��|�Fҭ��eh]}p��(��m�����W\&ŰĽ�)�V��Ƨ��q��8&2HR9��Gr@J6j9��1?��j>)�UtO�R��Y>XC�w9���fV���+;h�1��_q�#|��Ѡ-�~4*�v����M��	dP�5L]��h��Z��c�|G�BN��@��`/�f���_��b����r����i���s�u����`r�������)vH;�_�
��:V�3����^
h��v�l����4y����𩞛~ȿ�v�����e���YG3!�쯅\�n�|���m�QX�Q��8xl�d,|z���Rzp�a�#�� H��'�:h��y��D�T����<�!7G�`P�^>�85������EiNG�sF���W���^`��͖;q�ڭ�2�4�����@ ��X+�7�xz�ϑ�|�	�ؗ;�xa�qdiG@�p���n�s�sR��o���L�k��+�բ�ޢ&����FI�O�Q�n�R�P4��M<m�6�e���g2wH_Y�M-�̞�ß)�K>2K������E��LU�H��Qp�J�T@�"��
����y���C���!Q1'ph��G��fd"�uR8*����[�W� �7eP�P���_��t3^�}=��ED����{�����α��cS���W�a���TM-Z��j�^�F���l:�pݽ�u�h,�|M?Y�dh��K���$�0��_d
eNT��>���ҿ�CVB�Z�~�6�Oz�T�U>Mwsut���^;�����;��$�)��|�n���Me �*�h�k�s�+�J�������י�,���t�����<�����R���[&F�)c���P�F�x1hG��v�vV���V�-_���m�������<��4a�0�D�/��V�A�R�6�^xw`"��̘�����!o��x���DLT���_����V��틙{I^�Ȭ�Tm[�s|Qw�Y�3Y��I��|���u�9w>q\Z�œQ�H��9.,��O�Y1�U'�3����,��S�&�b5(-Z����|�7`���*L��A6{�QT�=����q��}qR;���i�{�]\�3]q���m�����p3\qj��w�\����I�\t��Q�ZX�PD��9�)���;�T0�2�&m{���oSP�*����I*�aD�ɺ��4\���܉��Ʃ�Q�w��E�A|�G����(8YC[��WZ_FC��㢼��u������J��Ѐ�J�������K��`������BbH� :�$4K�'��"p��\��K^F�R���:Q+��������I� 
^��a����0��Y��I�g��#
'��OTm���Db#�+��V �r׻��kcy�ı\����de�7��Ճ�)� ��*P��=��/щ1�&7TS�l�&������M~e��X�{ۧ�O�ۻ��1���w7#��]������(�yeg�}O�����̰)�]�࿹|��s)����A(�7w\�O���}���(ٓZ%��|%y��h��K�;�q���&Q��h
���=��>g���n�����;բx�J{�jn�,���Wg��3w�o O�`o����py&��;�����g��R �3#�[��e��K�5�!/����0�g���X�K�(4z�FB@t�P �5�D3�q�֡�Qd�����?2�T�GhvL��r"�@�kC_�U�6xz9GT�.�)�O�*|����m~���L�aѴ�S����΁���\����;����}�Y=>m��0������dm�����L!�Q�5���#h�.n �'%�4�k%��W��j@s����@[y��!�1˷��@�ϝ�Fҕ�=ߍ�||�l�CXPS�z���*��L���1�g��W�쓚��+L�E �w�O,�%N�L�r��m0z9�!�R��\G�O�d��l��u�zr\�̣)rS*�d뮭�`����p1(jde?�o��Ӛ��˩�c��7'ɔ���u&�."u�K&������Z�� {��?�W�������\}ڌh��H��!���9k��:{A�Q�`�5p�l���oQ"qʧg`w�@�nHL�mK(��k��KW�_��hD��/u%���� j��q\�m�U���J�b8���Z[����Ď����F�<E�ߪ�Z�W�����)
���?[,(��_�ޤl�^�vH�F�.#�@�L׶����T�$�7,!uC4�,w��6�z���׉�"2�"��]�߯)"I����1��<�*�p�付M�}|L�Ԋ?�*��,6��#�|`����zA���<�教�q��BUx;LI[����l�KX���K�K���=�^�%@�q>z`4����I���z��||��|��+���y�>��ԻC�)0_�pg7�a��f\n[��;@���� 
d�E"s02�-��6��pA�E��߹ay���B���2��_3���еI�r�]����.4[����mѣ���.4�M_�\m���d᲌\}��`NU�G���\,._���!m�`��I�x�-[���o:27�P+��-}#k��4(�.��R�E�J���TJ��I�:���c��]$�����!2џ�������t�($T�PH�-4S�L������ }��Sfљy��z�?�tD�V������YU]��p�6�k��T����* U}4^O�^H�0�̬Rq�/zS�/4s�&a�ѥ����^/|7�P��-��rƳ���9]�8V�t�����7c¹��UyE��� :qp��A�O3k	Ow/S�Z����r�2.�6�o��՟~(Z��/�'ʯ�����P��
&7 ��_Ձ{�F]z����װ5����N�C��Dy0	��\���9=����a��@�V��Z0�/��BS�k�@�������0��T����q�+��[��tA:9��W��P��U-����ݤ;R�$�"~2啡FW�r�o?��_
�AR]����!��捓	��Aלg�n�T��@8$<�`��]{�8��������V����m|�^1��6R��Q]1'�a`Q Î*��Oh���pQ�]��\)�V+}%-kkQb��Xاu������,_��x�z��ۆ;�|�����8|��Ϙ�V븸kR�����Eɉa�~O2�e�}�}��E��n��;P(vլ�g{2vԺ�ϑN.U܉R��
�|�"��B�r�\�1��⡲ʐ�R�ۡT���;h�5��"���o�ZN�g��.�B�zU*b�LN�RX"4�����N�́�y�ZY��WϨ��N� R� \֔>
1�w�n�����
8�k�/'td�9��Xld���$�|�,�Ə����� <�L0��'d0��C�7!��FYU��29m.y8BڕvpC������g�!�
�C��5�x	V��ڨgJ��k` rX;Su��<��@[uo웘�5�S�r��R�	և'��x{��W���s�E.(�X�t<l�a�Z[iB:w�[�uz����Ȟ�!�D�9pۧ�i2�O9��M��2�vS�R�;.�+��B;��Bά�"YEB�qK�N�
G���{�������a�
�p/�c>b�4f.��(~�S����t��%qԜ`D�x�fcqNڰ����Q�@ed�*i�k�9Ș��s�~��
)�����iݿ���׹��J�hU�rid3�ĬWd@h���ԛ	���s����#������p)��n�7����k�g�`�K�u��>ȷ`�,-�w\@7g�n`��{]k8��]��Q���S��!���W�	h�YL�n��
�^[��1�Ɵ�X!��k��&�N���)|��D���Al�K?��Y�t�?�
Rt���%�@���܃��Ss�y��⟷Ŝ$S?25f�P%�v�j���pF���\oh�-e�2�+Zz����xF���&+˜�vA�'������ ��Zs���'�*����~�$��p�P؃�°���i��uL�ւ�d��3�W,
[yID����'�z���4�`pmv)����@擮��Z^�� olH�P�.�����iy2#U�Ղ\�鱅
���}�	��<[Y��C�����W��i��F��Ze�\�C�,h�c����3=m�~?��c���L���I+T�pHdD�I�&�V�a�?�t3�̅ ֩5���\�c�V\Q���*V�GP@�#m���wcl�2���I��	" "� ���6$k��
C�Eu�γ'P+����i�"��bs�����S��墳\V��Dhن+x��CxW�
9*���68����������"�l�%��U�WԦ'lV%�pNxK��Ly�r^����rȧ~�O���%dr�Y|\�9�i���vyt�}$X�F\8ull���I� 2�����`%V�
?���δ�݀{n��e����)$w:"���ڇ���1��=�f��M^;y�ڭɫ��vF�{��m��[�#,��sPx�ZP���,�X����C��PA7�,h�d7⣶1q��ƜđX����2����B`�D���z=�dQ�UKGIC�쎳��WP�GA����Ec�bC[����_��:R�~���)6a=��R��9��R�7����W���AuM@O��J0�b�	LT�]�k��/����������<M����\QY���E��-J���c)�|��V���W����P��z�P$
k�,�[D3j�Ѩ}� ��fi����S��L����=H,���&����� ��� ��p�MQ�J�N��l65��@�p�A^.�b)_�6Z��8������8m���:� ]S	�������ƣ�c빡�}{�]Ć�n4ۊ`��.�w��S�G�Xxl)�.;�?d�����i�L��(a�Dp�qu�=*R���ې�Mc�gN�	��������|Ă�k5��K�+l�1�f�]_o7�a?wGy8���@��<ꨙ-T�2(I��sM@t)�T��QP�ʡ�UP�y�	�Iqc�i��K�����e�����l`����.wl�S1�2Þ�D~m�����:�&��P!��)�Ä?trw6i�����Lփ')T^��,m33�8L_�rc?<�H�w��*��:-+�vQ�qY+n���/u,�����P�QW�p��w�Ҹ�Od�@9x�f�G �k��x��1����4�N�Щ�K������+��*Ж��;̻:���_�1��c��!�:��e�|��6dM^99�����W�#+Z������7RZB����_f���u�0k�>�0d#���ރ��W�e�s����ǵ�a��FV��	{������_���}(h��0��+qŴ�ڤ���6�7��� �l�)0�2�ھ4?��
�Z�P�qդ�VV�׀yD���|w "@_�ך�Zy�鹝5�P���j,97����p9޶X�m�Ƒ\�-��P�����$M�n@���|�]v�[�%oki"I�wFZ�X�%D��O��Z5o `������2�Ѡd�>n���y�Վ=��M&����V�h�&,���Q����YhNDx˪uˠ�fU��MW�}�����,�MI��g�Ǒ��;D���&��bT�K��U!���\٬Bc{^����Ф�Ƨ���u��f��Dq�4��1������<�	�<Kq��3��ݥ���n1ߖw���P�s{��9%���:��xoW�W�1�������,m��8镒��2o
V��Z�ʩ6�WY�Qx��V(������ֈ�2}�^NB�c��fEe��v戰�sP������V"	m��Ҏ>�)���E��I��؆(�{�2|f_xz�}<㫷��8��q�5����b����] ��}$K�f��$���^q	��P��)������%���{�p����f%�7�[Gs��16Kߋ�w��M=&����S�O��ML����I4��fI���@����ߛM6�+M*�.�5�]����X���I�e��[�*b����1I��3���U�%����ddxy�=���K��O[��@l ���12J���<��U{�����n/}�=�{���~���)���S��N*�u�\�Q�����x̤��M�5����!z:V]������%�e����w�Y�K��q�v�At/���+���)��e�F0N��0^�<�W?O����9���f����A0M�@zxj��c�<[��r�D����TRB(���3�&���)I�N�}�I����$h4Ԩ�~��	��1����oۖ�In3O~ΉeQ���-��藍�O����@<&����@��wY22LL����UdԨ��!1�ivl�*Mba����BmȂ��.�%6v/���+:%Y���N2?3��gc_{�:陳�4�unfi:MR��]�<2�Y�<��A� ���+���6,���K��_�n0��:��a�F�zl�诟R�'
��iu�w����� �R2h�o�e���I�p�C�@�.��j9\~�	�+|uz��9�R�t�'���K++cM/П���α6�'|Er���Q,ո��7��C�������F�-��=�����+L;����L���4����)������LH(����YB�N�?�*�C���EnO��Y̡�Q�fϞ���j�������qt�{l�a���E�Z.���z�_��]�$DIvSP�B���K�F�������ö|	��}���f�1�Of����ii*�f�nj��Ia�Cn^m�A�!�%i#H���W9RX���K��пIz��7��#��p�$���%>�۳;���߂=� ��a�pH�'{�_r��b|Ѫ���4� J�Zb=���=S�@��_�r�Z�����sLw����t���m4��I�C�`6@m����3�}x���5�uH/v?�f�&7ߵ���<�y+��2H��x�����\��/���T˸�ȳ\s{������{j��<�A�#cڶ5���*y'�3T�y��}�n��P��R-��4�7t�Qmx3v�����5��M)��k�?J��~�ތīS�;кA񩎖Xdj��兊���#]˥.Җr���m����16�9h���������%�9�d� ���VP!���)LѥԭG���l�Q�un*���>�z����Lq_Ssw�čO[R�N�����I��	�p�w�	��)�����iy�<�q0�%�%�������XR����.Z$�����|���f�\�$g����f��Z?� TK5'eU�frB,���-���w"�m:=n�"��p��+����[_,�:���,6��*�l�n�g��wZ��������^6���p����&�B��G�I�o��?�Q�� ����]�E F�Զ$~�w-9u]�t�3I����^�/�+�i�]�����(�Ԍw���䥃uI�J�00��1�H��E�n���&̃����b9����e�%�I��׿�o�KXk#�(�^bh�ZDº��{ûfɤ��ޮ�zj�MC-X>a���]i�;f/0ꡤG�9G�E�{`d��`	/���+�1F�VDvrE�N�*����~z V�ܬ�Ğ�`��#�`�:��m�X���@Ĳr䤮����A�[��X�0���AkU���(0��a�c�3Yd\���fd-�6�K����{�&���=h>���_�_�2�X{1v[冷KC��Gt���9Qw�dHO��w乙 &��@�k��tp�+<�%��HzO�X4����{�py�q�K2gy��c��H�Rm�Z�_/��/��������k`����-�.H�w���í��`c��-�����ٍ����B�~�'��u�Y�e�we���l��c\��Nj�0q[l��h6��zI�.�!�j���%�3�4�؊?Kd�de���Y�['l,�s����<W��l=���C��īR��'��m�Ǩ�� l(��\/�G����Q+I�������Pը~u%�;�7���]��Xj�����o�lz;,��e�X�.�v�5`�%��}WB��E��0`.ky��vU=Q�~����M>De��q �Pݷ�/��/,�ճZ!��r��2ݱ'�i�>�x����a��P���$�7_-?�A������'q6���4B�=��o��K�J�p Æ2�6�o+�#2��0�=��諼�3ŝ��T�����`�`i{N��f݁cQG(�'lh*�N�"O@�Cx:�9�l�"�5Ә'?�)��~��&�Ơ�Ͷ����b�N�VeS�LrK�2��nm�}-����u�6o����~��݊��Olo�1i)��;gHs��B��6=[M�2��e��L~Ý�"�hކ�.�� y�a�;CL���g��z!p�8>B��� ��|�<�H 7���{���Wu*dGw�Y�}�E��톁�E��cn3�G�'-��2�o��:�L�g"ϼS���$%�?,�@�ӀR�c��-L�.�'dG����z:0M��0U��:*���
L���'��}�,{N*D^ގ��[��ҺF�&�	n��(B�8���^(D��?r�ψ�5��1� u z/�H�)P�B����m?��вH����8mJ�
^����- .x&�F �r���Oh�GM�L�pN���l�2<�W���O�'���9� �ZmZ��(AS�ۼ.F�fȪ�4q�Bt?���J�$�[�wc>�����gI�q�����*(9g��E^5�v@&.�[��������#}iqo5͔�.���Qs�k.�� �[d��?�9;���iߔ�}D��	ŭ�k�Zh�׭r�3V=i�BL�ф�k��o�v����+���P��Y=�}��M&��,��"t/��b�L:�<A��9.G�-]��Udpj�Eaގ>�k
=����&*w�#m��A|�U�R�ON�np�h���oA�a�{���_q~7�΃}�Vb�MG�)�:�f	a�/�Q�7�F/�.hb�z
J1"�@`�!$�z,p�a��p��>F�w5����s�X�i���K��*�7B/񂇮��?}Ԓ��@������R��T�����l���E���KF�[۷��R���%�N�����;I�����M~c�U'657_=�ŉ� 8$�!�:̄��ڲ_}Y�}��[����Y4���A�)�[��4�+$]����r���7���@�(�6���A����Ֆ#`p ����]�,�GMP"Y�>Ǻ�Lz'c��LGpt�F����J�p�$,R�u�ׅ0�N�Γ�B%:�x�>P�=�d��� �{��.��ZU��?PTP�0��!2��� +�׼@�L�G��:��y��,�r���G��JB@������:�g,�����fe<Z�vk�6g��B��
���.���:���&2��PV`�2��_��G�ș��T���f��kl�g�z��i�㻀Y9�� /�w���wY�55Sqg)z��d7����&~ۀ
0��4���{���� �p���d'#�g� �4�#�1��㩅��c��ewc0����h4[��B�s6�CZ�������/e#7�]���O�_2��2�ܤ�,�sz-��A���mv���І������N�2���+9h�6*�%;o2�2��S��0h=Yli)G�f�4[�$bބe�%=�hh�eH=�d~It�7���zM<Z��cLA��D���S�&���Q����>��z��+�c��w~A����d��� 7��.$�:��՛���w�cb��c*X�`�2�["����K�ig	���I)�3��9P{Å�d���#{��ߤ5EN(���Tؽ�hGq�h�G���D��x8�؟0��}֮f�y�r���z�������$(��M4�
�6��Ͷ�Ze�ɖ�t8�P��B��I����\2�I��g�ߛP�(E������ �dj�)]�����Q��p��Y��"f�l��y�D�*;�q��IY,u��Y�j=k}�[�+�<��hط@>y.��~:+�۹X�y"��*���y�Z�D�&g�V(�'�#l�!�}��y���Β��5\�g�2��c�����wh��W(hQH�"z�$YL�,繴.�Y����`�?(�`B��#8� �qL�E�����N��)�o��)=�z�:���H����w�������p��;#l�Ә�~�z7��_٬6$[��PQ�0��?��,�MiQ��O��l&DȀ����@S)�՗x�j�e,-�r��'��pC�zT!����k�^��a��E���+����̅�3�����UV7n#ē@!�7'�Ԙ�<�q�̀C�Wd`�J Bz������JW>?�?�	G5���<�.	��S����(���D�wRTE��d.8�t����챆��@�v#���R�]�z�D�_�^�s��G�f���A��>�D�lR���K�S�BJ��s�;��fC�L b� �n	�)�,�
����&3�68�����`%|�
�j׹�B|p6�˜vɱ�����3�դ�4K�L���f�#��D���E{5"PpӍ�#�=L�(���Y��ړ���CA�9û)��e�G@�=��sp�{5�V��N�U	���g���ks��Ak���O�:`�P![7TD�+
ӰT�y�p�^�E2��?
�af����)��. f+�fr�ň6��$ľp-���%yA!�#��$8���6n6'YH6���"\ˠ���c��r��s��ݕ$���X�r�c�V��$�or��w��ō=��>Ğ�a�;�⯪��`�UA0 �%|ss��%���[�����J�q�n6�S�Z�R�D��6�?��.�"�yX�(�,4I��O���,��~v����&=6@~P�{�b
I��O-pi��Ѐ�˳�oR�����}��#�}`tWL��l�,�]����Dhr��0��xbKٷ�{�Y���B����W c���1��$q⦰k2�����e���{��ݵ�C���K����g�x:���pv<���G�9�d�O��PPy�.���H�0��j��2;�Ϟq(�)����N/'��}GW���e������7�����ɝL���Myw¼���M[K�}��9�rԣsRl�;�o9�861k2���E����'#q����;)��#����RN��0��9�\�{Dpx����dZc�����J5��RiE�����W
�6@ƃO��]Z�%e��^��tb�	�f�oNT~)_$X�`�a>V���.��ʟ��]]����~�_�ǔ�h ��y��/�}��E?�9�@�*�����A/�^�\�f)�Bn����|����̧�A8}����1��b"<�R��g7#���8�V�߄�y��dJH~Z]W�e�c~Ѥ[���)�w&L0�~�D�SV�\U�Ǘ�u��(]�H����fĉ��[41h6�ԃ�BW�έ(\z -���/�:���Č"�(�C��<���$Y(��~Ͳ��{�Dy�C-ki�P��
��O�/F[�sC1=��ж�ۮ��:5�)h�>Ǘ�U��p�	j��vЧ�E�ַws[��ã���³�qЩ��b�mj�gr�W\Zt�g�������H:趫��{rn�n�_������uoI�d�`�gc�5wQnW�r�x��j��?�9���FG��>���u"�C��Ⓢ�տ�EERњ�ᡬDL\s/��{jօ�R����_)�˱Կ�I���ЃK���$�������lMu$�6ոd����l3���d�w)�?}"�it�(�Ҩ2A��0���u	Ĉ�B�Ιj�n�")V���ڞ�Gl��eZ&�犩�r���A�k�{XJ?�IA��9���(l�|�*`"��\*����aި���>�aC~b!Z����h٪)��p�e�sy���j�_Q�zF��Q���<�T�>,�V�G�/1�n����m�<I��@.c�uxn�3��k��,.Xn��<@E>����}M��m��*�Ecβ��r!�S�NG p�ۀQH��c��mZ@��0Ӓj�^�����	�Or�xz��Բ���*8��Ou���~�q8�Ye}&`_�j�f�~"-�ۊ�� �2j���a�0����s�PAU03LBK�mt�Ɨ>V�wӡ"$O6t�݂���g���׭f<�7��Ȯ�K�h�����`{��~_눉�\ T�_<��x��}[�����h�VY'��>��CV߾��0z�#�j��3�0��e�1Ҡ���{ ��w��ߚ9�tf����d��

Ӳ�^	_f8�9�n\���o ؛�/"�$<m����3���7~��y���lQ�����������7�}σ��cq`c�uD���M�g�vs�Rh� }z�F�]�BeB�l~��@ɒ��j5�/P#�ٕ��_����v�;Wǂ+Ğ�NW�G���=��7�t�����>o�>@�xoL��RNG��m�WA�K�P����}I96Eb�S6`GLǖK
��\w%�l�yg'�8=C�[B��G�CblC`J���]��/gP���1PvW��N�Q�|���@������-���:+'�cY8/��;��,`��諏v�.���!�}`7��[t��;`'��F�y�(���K��FK%�ks4�Q_�^�W>�������Ѡ�'��������_��Z��>�Z��R�+ӯ�����Y��j��6��X7�g�r�@�� '�3/4�.����ó\��*-����v��}�=���?�
��Iy�'���� ��0���������n�ya���(P����L���Q
9�8x��9��(��i�T�@����!���0��#��o��g$,g���ՋBƅ�� �2�0���LKͤ��ݵ�������E)�H∩{g�	K�d��S�3�]Y&%�����|bG/t/�/�Ȼ��5>L����W_�,��NڴW}���� ��q[�>GgxY��{=]Rh��7�ލ�s[��s]��Ѽ�6o2X�'���{�hÃ�!jG�=GzA��~���J�0��q9d�-�9�-:�����j'S ��"�&[r�O��d���*�-���c��_Ɛ@6}���dQ�=��5�u�á �!��o��L��:��&��[6������D�Ӊ��O����H�)���}�1lB��
��-��$P����ޕ�%�����R�cC�.�$0�F��\���������-�a���K�h��t�7�t�*�i�0�0P��;L`��R𿷤8��Ϥ��:>����{�O&����[��Ά�V�F��G��U�h��\��s ������GLu?���\ �s��v�\���]>���Zkd�A��|�~�Q�BNO�y�؞�Y�ݹ�=dพ��@8S�n\(���]B5������{�
A�E�ziQ|��[6����W��|!�Qs��H[�=�����A#�}Bnι�٩	'�k�Y�Օ~�C��ݱ���`̏e���}��X��r�/	��
y���4W�Hu�~���C%������9��3����^�4^'A�,�9�����AsZ#�VY��9�FQ�$?C�-]b��C��͝>A���-�:4���u)|i
t�uuN�,R@� ���&��p��Bp����5���t��j1^s�6�A�L��4�gC�g�_������L�p��j���h��Q��M`��p��iB[�O\�1��NB���;i�~N 
�Ɏ�����7yK���Q��Y�r7��<�?�48򎟺Z��\5tb�i�Z�8'���sH&|ɄSiTǇ"?� �ws:��ewn�,n8x���:�KS�f��^� �x�tH�� �Q} I��o��=�wdm�Z��y�k���Tv�Vm�\�^�&׋�MVgc#K=W*���jQ�c1%�� �V6U�u��cy��p��dl�z�C!n��T 3(�(�u�%ЁnQ�c9��$C`˕/�����	�
� ;Y=fD6~o�	��k�f�7������ pf�/F�.>*q�*��S��;5g��\�6k��K��i5����؜W8�ɀ��B��5nSӫK��dI!��d�:���*4~����m4�m	���U���p�G�¶�}"���ݱ������MM���2�H)o]��S��O!���P� ��n�>O4R�T���௥r�gk�k.Is��yB�ŎAM�> /��~�6�+�f�L_{p롦��|���GPFH��Q�u608���'tKgIg5XZ	��e>�m����?�\t�JnSJai�����J��	_n�}L�Y����^z�z*�keo��fc�^�nQ�u1�#B���pK��H�'poDQL�������M�<T1��,}8���fd�ӥ��޽��>[�N�ˉl�[/�\i@�e�F�[���jpD)gtYԃ?_�:��A1�����LH�$������z���s�Gf=਩8�V�c�e����cR��v���.׬���͂4��p�N_�C`�0�[��#an�-��@�$�Go����'K1�6-9#������»��}:�7=Dz�_7IW�ދa&�p�Q��>0~E�ev�]T�>�$`���G����"�c��
\{b q�m�H�(枮 n�ē��@�-5�1n�W֝.�k���ɳ���{#��'Ɋ��/a. ź��(�q�ɔ^R���7��W}�r�Z�F�A��	7���3���ޘ����.�b���U]P����ę�Q��]���.˞{n̄g�� �`��vZC9�(A�\���$\�%��s����	虿�Li����"�7)��l6��I��f5��o8��h��LG�݈�T�)�>��C^�W�Y�ux��J�zF�t���5!��Z���/^rEE�>m�HkF�E��4�V���r����
;���C������4�uY�gk��c���Xb^�$�{�Csܟ��嬹{�	K�I�k�B!���W�Jh�d����[�wB¥[�����4��#�1�4&Z4����Ɣ5�.�H�¼Vf[��?\Ƿ6	��#jϚ����Z ~�3l�
{�Vvwx_��ѯv��[v*����:�A���8\���X��4꠪� ���Y|2��a��w1��ܓ0��n����e�m����:{I��7�]B�w�o�����1U4���d��U�м��ң�}����I[���Զ����ˍ �,~)1���AP*�5s��0�ū��j�<�����ߠ's~~s֡����6� ���s̏����嗨�'@���/��J�A�: ��I��YQ6g��yv�3�E������� d��f��R��L�H�1�;l�(Ro�Cb2)�Axb��J�ط����&�k[�2w�3g�xޟ���a����!niq�u-�q$ΟK_�L/ ~K�gvƬJ�?R]�]����D�עR=X}��/۰�`���.��B��C�K��}���m̋Vb
�1F��!��x���s2`�/t�Ur%�����]4�aO�C@��Dd=�Kn�ԭ�ҁ��� ��(�>EƱ ��?f�#�J��mb�&3t���^���9��z�h
N�94��1th9�k�{��0c�xh�1��H�����(LGR>���9�oG�b�s���(q���{��~˗�f�m�B~"�W�sʉ��-�Mل�I�;Y)ff�ł= ̺]�a���"�T�6�&�O��[�Y�*ei���vի i8�.D$T �,BL�^����_����2 �x�-��*0�c-C�y���l�9Per��B��qU��S�%�+��;�`d;p�ϰ/�'=(�&8��A+��Ke�h������¢n�륥�,��.h�7�w1\���L$)�u�~���ME�hԄd���)�I��W��s�h�NB���zn��wN���V�?�����!�Hgi�+�̫1u���}ߜ���CO�g[
��0��&TG�C�1��6�DcY��!�a$����씕�ڥ�y�tX��8���o�Z�K�"��{*�z'���?�\x�'�A�K3x�O�*����b�R�'ц V��GҪ��?������m��L.6���$�tx
��~�qb��ؼ��v6\�H�̱D�,~	����� �2����Jz���U����k�WV�Y�V$�f�SS�\�/,��v&e�\M��a���2n A��m��I�'R�m�s`��`�����
SZ5����-���
H|�)fp����$����t�Q�z?���?|�{o����&ˑd5�?/�v�j2m�7�"ņ��u�_�; ��g�[�c�F���>�g�e���Ѳ�sǪ悲1^J���ӳ�$Ϳ\	�)���`���]P�9މV�D����L�r�x��r	s)x���mg�s�@A/�� 59c�#_Hm�߷���J�ҺH�*N11Ж�(�/�@!g�0o�����g�3���^k͐��Rqytë��>�Z�T>vmk$�2#�Ǒ���O�0�d��:���8��p,�Y�r5�E��U�f��sω ��XH>Ѓ��C�9n��OKDS��u��U
fS<J������v��ݨЧ�wW�c�x���`��B\�v��� P��O�&��eAa���De`���P"<�lvX#�r�h[B�7�P�]��z�{O�D$}FJ,n�}M���䷤�ܖV�������2� HV��]q��\���Ó͚�g&��Ć�nx��C��� '��!�Na-�QP�
���%�3���v}��s��r�k�V�zp�Z��BSg<	�_*
�Ȏn����"�!y%C�-��q%���P���2Q�����j]�*%m��VIoB�}뮷�����w�T@B ۓ�?��V�:�I�QHk��\j�m��M���[Ò�i��4�3�#v��6����j���
y���������%dH؏؏� vX P�����¿m�J��Cj3t�`"j<���rd@=Ĵ&ӛ�q�~�mՁB��۹�vې�ga�#K��#�����e��>��EXk��G��( ���0�*�E��Lbj�o�3�V��WEZw�����b'�0�">�ʚ:D�[5?#$�p�g���Yܖ��>�<,-*m�������\���O��Q��K^@_ꁁ��l�� �I�����V殘�����t��lN�v^ �!�'L�2�1�|6{)m̞����C������;?�}[K��yΊM̩(��4�
27��4�8؀�U���&���1���������m�jri�I�k������^1�g'b�ϑ��6u���(	�J��!���t���I�J�2��D����	�h{��7�P'T�T���q�>�M��*p0˯0���+�G��'#��&�K:�PL>W�S���@X>I-x�A
IAx�Td�b�]�=��&ۼ�f$�`���8c���Ž�����;�#�/�~�f~0���`#�762g����	�3k-�~��j��"�Q�M����ON����0S�R4��(p=��܁Dx
q�����[�s �I����A>��Vt��e3�U����O�S:��(�z��ܛ� ���R[{��E3�AJcI?ҙ�U���>X*���ɜ�{pI�/��{�7�Ae<�nulq�b9��::`��� �5m�"�SI]]�~����c�����,V�:ma��]��!"75��v"�C��o��O�
HP9ُ"�c���,��ć�iA�U����np�^�[��_�\��b�?Iv�=��`�b,(M���IDˮF�W �Q��F�(�ۭkZ�Th����U���(t��̨q*�}��\դ�wL$#�д��3i��B{5yBشl���5�ͬ�?�؁��Y����AjV�"���g�W������_j��Me��٦|lK^�ZU]v��xa��%� ����<��=��7���-qΠ�<���n��5��%�|�ŭ��@>�P�pɐ�(wO����$
�.��n�*���}�i�$�?��8� `O�Q�aG"L@�0H21����bs#صc�(C�@��]�͕��B-�E��/����H{V9�f�����z�X�Iψ���2V�ɮ�)2���g����b[=�o~�s�Ѻ	zf%���$��Ԣ@�NZ;T���JQ��aT*J���S>;���T�N̋{�"�5fI�������ZQ����An�J�����r����(��L�F�{���T����H��e����RjMF�H�😴$΄��&-;^&p�/�O�R�l./ޕ��A{�!e����!{p�[k`��Jb��+C���U/�,�'D=�sk��6�	R7�_5z� ���"ġ�	��}A���70"A7���\,�D�mRd"�>��,\s"��o��+&���(M\��ؐ�$@��x�RDds���5�����>'<���
sz�)m�ȋF�q:D���q���̴�k�ph�]��g�.wY2�T>^O+���-�1.�o�֍C��i�w��s;/`�8����N��v����\o
�O�b��
L5��l�� �{k��������b�c�l�C���x.帐�@��h��#�9�ИX
8'�\�UP�	�&o8����y���E\�b�nZi�X�~�I5��0�� N�EwĚVMΊ�-�������e�D�}n�~eLZ��r�z@�H,2��Gj&n^�	�|�n�		M�9r9>/B�*/"3o��(�c�\H����q�FF4D�_E�W\0��B�q�qq_G)�4瘴�xz/˂xW �D��4ZWmމ8Mf�����L��^�ŢB�c�Ț����@�V������lԐ���^Z?g�<�f���$�ɸVG�E���p�W���"��%y{a�rkh� !t�UDM��o��\��y�u�!�{�$��c:�2�I��J���J�"��Ni���]��:�Z�R�e)����ӣ������q�1��
�e�ɸ)Dϗ0i�w�J��n��G���� Io��sʹbZ��(#��O��&U�1�;Ćxq�u��K��#+
'�գ����(�%�7��uw��~cO�(<2F�G�\���)i7�}�%�������>K6�~x�q�<3*��_��{�]n�_�c��YZ�-��c�;��39��ws{#٪"������9O	>䖈u|����"߷�OKh)4�e)7��<b�I�<(�m�0��<f��	Ab,��;����t=0�<R�4�`xf�_������]���h-�qPA�(�T�Wi�N�#���e��z�JN���L��T]A([��!8Ey�tVp.͝�3/y�
��O����8���W��PG):y�U�H�g��ܮ�7�K]�7c�A���	�,Gx�w������a7['Ϥa t>&�����SQ�b�$v�h�t�SxѰ	t���6��=u�!��o�2�a7�� +�v'�Ypc*��,����10T�_z�(��ǾR��
��	Kk�F���v�X�dgE�ʏ����X߼zo��u.b���Q�z�1fe�Uid�&(��,'���0�wӽV�1�N�Ip�Z���t(m��T�;زmb�?q��k�O@s�ЀΨ{L�\�UT!�u*�����mR���(!����Jub��ud����ۚ�@���r%����_�R���E�	A��IP���i��|�3|7�	Ĩ63_���Ҩ�	ea�t��.��=舺��f
E����ډjc��K2�vw�.U�Q׼�'s����I��*�ǩ�C \,���7(�v���7�.:1�1����vL^�-$��Ҩv����e-"�(5kFQ�P�׽�@[�ete�*�ܽ���w���L}S'*ȃ���c_�g������އ���C�#���6�l�PW�,�9]'�n�D��t�_KJ�PE�r�����9=G�6�4�5��+��Y--_���W-�B̲�\��u8[j�,]$�	[��U��2T���)a�a�A�V�#C���h[�#Z�����|�v��i;o�%���S���9��Z�x��l�ֻ��+k�G�{8p�u�anґ�W���P�&>���53Y�u��F�C�e���a6�iO�FǐU|m��s|אM� ?���6��02�Qyx�*��hn���{��Ĝ+b��7n��y�N�3U���P�imc�n���{孇��ׅ�8��	Z"dU�8������Aj=O	�F�O�V(�||������ϭ�2�A�����)�/"�-�T�g.tSȓ <�rTl�W���L��汆58���~�.<��2���~��<�]��]�aH�񔼤�`���0mFJe�;�ß���JTB=�W
��<�O8�YL+m�P�E�ц�<FE諦�{���lO�Vf�����0hG�(��+i+mt !$k�Z 6m�#&(.�x̰��k���/�� %����I�7�6G��)!)��
`���뫀���Ց�dv����%���iV2Jaa������6�I����T
ާu��Oz�c�t�_+30�����9O�L�!��Rq%$�Й�1BM8LghH�83�<���s��{��N����j!�<y��h<���(��-�ilix��\[ؗ#�/-Q�5�?�
�!��-���E��i>*ΙÊ:B�(-�7�@�6�A��T{">�Y~1]Rw�ˏ�@��ɿ�[el�q����Z�8�E��zPw��#.(�ʣ,%t�Nɜ�؋��;nu6>/�k+R��PJ��}IÎ��`�F��jf�H����nKx��|)��x�j+c"Wa�BE>�%9�k2p��#S����,��9P����Ң�,�nW4Ű�7��A���q�� ��r2����,Y�^8���㬼v���u�5}�Q��d�0����g��qL(��h�T:��NB>����:=�l����p�M1r\�=�0{{K�7k�F.�B�[����B�%qǽ��=L�M�;_�sM��G&@xN!��n�B2f��L�/�(�R�y������_��3:DwJ�5"���Bײ�oԭdۑ|�B/�s��޸���B��:;��E!���6^RHf0!D�*I|ھ�)Z���؍�� I��*���X����?�B}x��Z�9�}�gZ10iR��P#|e�:�.�?T�e�?j1Tћ��7�x�0:E�vP$�M|�ŧj,~��Z��,��|}�8X�߫�
��x�&W�^��
����~�L%��hjV��y����k���Ӟ�A�?e��gH��Ǖ�������������$���z{����h�??W�Z�����Y`jThzn(�I�.A������ی�$�}���ڝ��٤�8e�~���cDvd����-�WV7=�|Î�4r�����̕1���;8?���y,�Kʎ���'z��5>� ��ʮ�w�䓲)�z��b�PPF��b}5[�-����!l0w�4X���\��i�+��ڟ�/��΃f�nP:��֓e��+����.2����/�؉_]�K���Ow���CӀ��N���=�$Y��*��mѠ�M�u���\8�Q.�т<+������0bus�������\�`ȳ�ΨU���~��Oƚ���D\�]G8y�2O�y��:�_x�:s��;C��q7a�|:nme�yD�ᛠd���ao�O�]P�*�Ϫ���oL�|�؃��c��mn�Rf�(�0��ʨ�m��?�ժ-��Z`<�``�x��D�yy��⇧!�po[V��\�n�/���sg�ܸH�g���	�k���g�}��K���1�����s�D 9N�O��dPv��W�i�t��)�v�Q��q3ħ?�b������֨!�;?%�l�����)i�!�IrXT�Emd3�sMoYV<�>�:b�Dz%�&��Wӈ�-�4�M���$�W�
^��&��H�%��B�`F30���^�_��u�t�M���?����Q#wR���f�����-�O�%��t�<���jt�XT�]}m���cphz+ �@���F�L���ê��.��	�� )x�,X5G��in�@�{��ʩ��u���Q����G��*mM�����V�e�%0�3�Ů/����
�낱9��Lp����h���s�ZH����O�������)ª]�;�@Q��3�G*��N,�3:�� w�H�>K�-�h4����4� ^hl�X.A�X���iQx���-���/-���08�7I��os��������J�dLvU5�v��n�����з&�
t�<�&a���&5� ��1����$�,�=��{�� 2"ʙ�]tN`��\k�.�LIt��x�@�ɹ���f��3�l�_g�-���HE#>ں�¬)��{>�ҖO7�W?y��YǈL��Mŗ��f1U��uG�+R���x{	��f�lp�����wQ��I�7�Y��1)��e��(���S�&��p#��s9�}��	6�ɛiW`Q�/�FS��f^X
�5F�aZ��B� �(R��2�M���#�>��?��0|��n����}u�SJO���[5��8q�EQ�%��"���<A�H+~�M��O��(��?�;nUg�lV�Q�)|��_�04��n
��e+Դ|s ��_5�`�r��G�Rθ�M��"Vt����$|��AU�,���\yMy���ś8�9A� ��_�/x�����/g�5�i$����I!�IK��?*�����*o�ȫ�(�S�����0�TqKϯ�2����H��d^N|_�vg'��K�k�ĕ)2���W�}΢i���.��?��x�����<t���,�s��av��r��'y�&�g�^����;��������H�8�W/�#��6z��3dfg㜤�Cʶ��}��
�F.�-javZ'kH���Z�_�ՠ|y���Sl'W-��E6���έ`L��T'�߯���[2(ЈZu[�ok�J!�m.Ļ���"a��f_5{�C9p��X}d��1��O����Mw8ҵ`��#zf�FGe�X����G֘N���&[@-����>d6�}�9�j�u8[,���n�`h9�����%��x}&�Q�9��ԭ	b��'�z��ѫq������Q���4lp76�������������6���&*/g�mU�g/Z*�4
x�������<`���R�F���YC0�#�w���Qn&P�	�bN$�+��b|�Rˍb4~�D��+���d��2W��n�+�ȹy_pؚ��dc)<ﺵ
����>��묜�lT�6̤ފ�Gli	�&�ڇ?��w0��?�e���/
]�f�x^�(?v=l��P�tDFz���DK��e<�x_��	�~fd/�SՏ��`P��,���[�����B(�Y��b����1�G�`
^ȶ5���X����Sc�Rr�v�sEA+�\�{���=a�{�JW0v�xXH�4ݭnsϛ%`��c�e�,,�:�}��o_��𫔇�/�ch����a��QAC�fW��6�N�y���q����S>�����:�F�RRt� ���R�f��l�7����_�����������#Y�D�`&���bޤ#��7vC�}��r����r���P�$4F.Y������ӸW��m�<
�/WIܜ�Q�ǚ�D�a� E�?�s�(�&�<��=s�:��߯�H��Ike��H����˩Xڐ��L���M�O�HX!-k��ˉ���^tQ��.�"�[H�KQH��R�����y%���y�C�+NpS���ӥ&�{�/$�L��8% ����YaQ*��L+�����6c嫄� ���{Z��?�x��%��.�
m��'1�p?dL�U7tjuf��Wm_.���%�n�&��6c�j"3�0
Hi� �-��,m5�c�P�'�#s5�\���S\�-M�M8� �g��l$ �H\��b�T���y�>��t��-�x�����jD�v�#��ߦN����K��n}�<��}*�ƪqB0L��D#X��0���������
U1��H�����G�9>R"pjt8ف�z�m �i����<Aܙs\�"�F���ɉ��y����U��/��.��*_��ꞏ0�����|"V���h����%�߶'����ײ��=oP׌��]��ػ��Vb7[c�K�I��zH�u�Ǩ"��s��w���������p��soC��xi/0q��ϱ��êX3/@zq�`|c��
e�&��u�ŌnkIƢ���%�이%Ò�m��w�)��������Sc�}���C���	�Vr�/����P�1�Z����Q���t#Eᇼt��è���@�ZH¤q�LTE��F;x�FOQ����Gm�O���g˙O����Ѭ���5�+���!��������ۻ���m/��<��d�^���7N�h�d��jT���NXz�GHqΑE-�ʽq*4�9�:�P������4;�����Q~�-�f��'Rll�U%I���N�C�p��')����:F2�뫆ᇾ2��×r�r]�<b��H����械�3�v��n�VL����(7�±P���(LCD�.="%`:�ݫ���MJ~2F[�H^M6�B$�"A?�Z��/6ߛh�!�J-�`�X`�0�9ٖ�e�
6���dǇ-��{�Ȗh�ac/�b�7���$�ݠ��^]��}�g�m8^~�:���pgv�4�͋��d��
&cd�|zR��c�F(��_�0 #�e�߁��%P�E����|k�J����ۘݻ��L ]���V�rf���U�z/M�|~���)4�I�꘸i��M�γ�a�Y���DX����!������.��;C����\����"��`���m�紻�Fx�����3G�;�p��x��F�0{�0IeЈ�X+sxc�?��/��O���aLx��n�w_c��p1�ɳ��a��DŘ�)y��������x���P����	�XSf֫b52��7
��d���;<���w�Y��C��[h�����#�k����i��' i�-��G3���2�W�1�^�'��O4�]Rt�}V�mux9�ړ���pR֫\�'�oS� �ER�^�ck"���i$�(���o}��52O�t��ؔ'�V�|��q曪[߯�>��r
F��IG��a[�Q�!���Tj�O�&$E�Wmw<��AdլA�
Gq��V�-��m��`Ɣ���U��Kqr�,i7� ]�!U��������gl�T�'Q`�ʼe^���`�/�wkI�}��b���N� ܊���L��羅�X�D�������7��<���:��gitl�n�Ư����FdVocQ�O�$����4��E�y�����ʐ�N��O��8�c��1#��W�K�Ļ���sb���!5���q\#�C��ɜ��jF��(���K_V���|�/�3�]����eA]�>L�T�n�r��=�,��<~.$A���V�����#����-��>Sa�%��G� d�?X�3��s�������)�j;���
;�Mʑ፹,��uL��|yvwHf>߳�UZ�����O�:e��T��~$�92���'T�i�fS����k�O�ӻ��+�i�����Z-}t߫���ڥ��حsh��|n������y2��+#�-(V�uvf��D�(*8Lrt���}�$�z�	\,�śv����kH�X�n�a��J}^_�W�[V�ͭˍ�#�L�פ��s�䃦���a9�{�땙:���#�4<yg��D�3|`�f��7��v"�I?�ͩtI�^Sm��WJls-�q���i��Sde�����l�i�ˢlKd�6�WJiq�[����-��h%+!�4�G�L{��fX��-I+�&��� 
NMaO��<�b6+�F�1�b ��������1q$��iƬ0�H���Е��`_v��tpo�?xn�7Ej��K�Q��vs
�<�p@�L)�tθ��vFDو�<L��g�$��S9���V��s�� d�m����̂�0Y!�Q�Ӽ�I.Z�\���kʲ�@$�|���DR� �#\7`����ӕ��HXh�΋���C�\���d잷���pت��wit�o=4�t�����5����M�@�ߊ�L����CB�D&1=k�g>LlMc��I�����ID��"��lz޶}ړo���/���[zR�~!Qk!;_l��[ᣚ��Cι�z^4��*N"�W�k�7���L��8����Ɖ��7�.�άWy-WY#B���V���"�`��w��d��k>h�.��,L�A��&ӖގB�8>�e�R��h�߻$,%�z�~�~kC���~Ay��X��@��N7��l`(�'GS�8�2a�̧n=��3��jZ�HTU8�� �ǲ�k�:}Dr0�]ձm|ng�ki���N����Pq��vm�����o�:8?�-���hj��F�qG���^ ��V��������׆�=zkWM��.�Z>8?�^��ۧN�A@�j�V�D�J{V J<�L��nCG��C����[��O��+BB\Cٳ���ӿ�)�H-vx�Jؠ0��f����8�f�z�?*FkW{���&K׻��zr.#�~�&��o*���4e���B.�?v�+
ZȾ�C�V]�G�<���uEr�ez�x#�;n��Щ�^��WR���꒱V�����ӽ���/o9jy�w?n�[\*��`r��pW�H0��G�bd���u`jn;�Z��HC��t�'4$s��.�k��� yq�<�$U��M��޲�%��n������բ0ې�Ioխ&�<��c`��Ħw:y$ɑ�3*5�\�����u���j�̽%���Vg��|�L)Է�aq�",����"y?���^D�τw�Ci��kq)�B�Bq	���gf/����ʬ���(��z�����G�_�������`�*�Xe��-|:�L~�	�>��n����sx\�|G�ܜɡ@-�����T��טl2��k+{BzZӷ�ʝC��ۊt���)��ȥ�a�yX�U]$�|����n��iYvД7���\�q�7ݳ�^��8��J����]tj��g��|�;T��ڒH.���]qo����B.K)�[L�ث��E��ErY d�yL��2Z7�yHP�4����O�d7���C!q���d��ŏ΃�} �	�#����^�ѧ����1)�w� ��n� =�!T�8����ñ8t��Ћ����N\O�=�l7 �(���"�6L��ye��v��:��A�� �-�j=�R����{�:N$����oJ~�g��'PE���I��\�����4k���G8S�X��4$Z�§֙�t���ƈϙᩍH�.Gm�� �v0]��ɬn[XE /��{��3��L��]b{Tr{�^�M|�!�a������r�Q�I���>�>s��b$�����/*�H�hv��+R�f�L���;cu��,��i:�H���[�=Cw�%
/�ˌ�iOx�w&�N�]p�_9TT����b�p�?��ؙj�B�:)��>r��jVo��8*X�5�պ��?���{*"pp˳���lN9w"�nu]�&�"6*-�I��X�a���ytQ�6��D=��.}�����QS�CQ��H:Oɝ���X��x�Ҡ�F5�;*%g�P��"9"��ln��ڣ���>��~�U��O���r/ު�ǥ(��_>�N@^dɭd�)W��+9�[�����~N���pc���LւcU`���v�w�ԧ���ݞw��]+����1�Ko�^������>�ԃ6.oǵ�<I�U<Z��V�(�$S��Ezj>�q1��(7��*:~��7Ҧ֭-ܫ�łV�!�`��❧
6�{�����|<�=�.)jx86{�P5[3�V���>�5�O+���WF�S�l4�VJND�c&<%�;e��a5I�*����$]��Zu����]�1'�S���|޴�y�t�G
l���8i	>"�D"��$.�<l�� c��%��@#��?�q�Q�� ����A:# �:��v��ri��̟�=k8I�?'�'^aV��12�c����ڃ���lոN� ]r�F�?���r���`�K��W�/�ܺ�(�ijyV��~��G�Q������l�������P� 9�m�}��кQ��W$�۵�V�E����߼�����!�YXրȔ�ǚ`ؾl�0���ÜgZ�����PŮ�h�r���֋��J��E���a��S�E��Gb��n�R���?G ��R�W2��0w�eC��Φ�(��L;gï�O�vv� �����x�m�8&���3�`-b@1�����SV���D$;��� �@5�.� $��h�
<����D���r�� �P���#Pg�Ȩ�E��Z��Z6%��,��m�7��b�R]};�A�&w|��Z	�nKڸ�����ʗՕ�|���-oJ�a�2��bK���E�ER��/@� _�&{iQ�ó��)rь��D��fc$�^�9�C�����rջ��)~e��<C7ޞ�cة�t�:��D,ٜͺI"�s�ù���ڍ��q93Ѡ.~�~�� b��|�J,E;I�tB�k.ǓY/��^XkKBԏM��N	�5X��7/���@�
�E�. �NM=!��@ix�Ir1�9����7�^g�Qh7Ə3�
|۾�@L�*k�I���;�Sۍ$T�okCm�]�џ^&��ta9��#�X�����)��s��N~��|@�
p4I&�&M𱿺'e/����$@5��It&H���(���xA�������E�����/��-����> 7�ɴN���>�P�S��ME�sP�:�$���M �E۲{_o�CM(��&I����h���5��`�B��%,�Lb����Я�8(�������)C��y2���)��ÿ��P3��íA/QJ�|&/��m����<�Ht���[� �Ѫk~��R��z��6�@�
oM�{o�| ��J0�(��b���r`u�M�6[�����i_�0:|8+��a���N�0�2�o��e�)F�m��� x�|�*��g��J2tURO��?��:����D�����r�LF�om���[�t!}(rYb4��ao�΅�.Š��k��ɢ�u�_x���<�̨�9`�p>\�/�ȷ�a����_j#�� ��F��:a��2��G�����b���]nWoG�b35[�/͵����.eO3澕���H4w�&���j	SԣP���D�]p�2^���D�Ek�a&��@��M��Q���r<ƻ�|� F謽��z>2�}9�躌���ͥq���kQ��H*�]���ο�����:v�h�� ����� !fFxX���-ŵ&,���v��L9�~��(�ͯ�s��9�>�T�����X�|�F���J�"��L�羕�>��������?2x�Y��r�f�" �PbE�g���+fMԗ����\�	W��Ϯ��*��{��'��1$)�k(�v*��2+��$z�L�Xf��X5W	*��]�����b�+�N��(�����*Q�P�ѣ���������ɦ�-<"��A$����s��Ԧx�27�w.���%	yP�����4 ��I�?ɤ�޽ppK�F|]�
�k�eC��?�߻+�(��"�Nڟ��mA3إ|�FQ=��'3[�o)�0�)��ؖ���ō�?8n ��ύ$�np���*7����Ŗ�כVa7�C0-�ɔ=��� ��D�Vaߕ�|f��C���R�
{Em���Jj�. F�/=��4��ع�+�Oh��#o�-kW��n��y����/�o6�����v�.����Gbe��^��)��2�����oF�$������`�6���ʌD��圗��6a� FP�p��Vx��_��uTNV�ޞZ��	���]���p8뼾�Xµ��t�<ºݜ`�ѵi>nP��j]��
?����ŹN�.�Ch&h���׸0���gi���i�H��A05�ͳ<�%�TP�i^7 }R��k�w�~LB�ޛҕ@��҅�6�tL�C];�̯9���7k+ �L��G3#�\��_\��}!]Д�'1�|=4�_�鈞?��J!3F���Oq�'֧[ަ"�3,(��F�q0ʯPQ�����i�R�H�uE�3J�$^����1���G�rGx��E�3q��y�`���;Z���_�K���T��`��΋�7:rG~7��<%Yk�ܒ�+�eK�(��RTw�P�
�	e\��4�c뽝�%f�K��PPr(S7RORm�Z�Rm��o�ֲL�y��_�������b(�cYS:�)����0:.�)��`�>�,K$6aD;�[�~�<�
���-i����mo��|#�I>�xV����ߐ�Y���$�;#��_��+�LQ(���"�n^�G��(����82�b�<h%��ݔ����h�}G^*���U�I�?U7��zԊ��h��Ȑ,đ���Iw�\~�9_ ��V�ؽ�o\��3�}�٫����kE�o%X��"�\m�!l���ۦ�񠤉�g��\/��-�k��=�,~����@���Ԫi�$�=���~G#��y�)�%�T�覽K�wN�с�� �S<���c�!�
�5�Z�h
�풓T��}�%���J�z
DÙ�z�4M�ѣ+1!����]��:�5G��4h}�;9|�J�p�Mz�%�M���S�?c-�u�DhA�T渼����fB�;<�;�3�z�{�M�ol5���`::�G�	\�8�pn:�p��Q�w��!GaQ%��ttY���m��芆e�fx�#��x�1�U����=}��i�����/�(	Q�ޛe�i07i��Ԓ+V:�諿�nQ��/�>ӜJ��5��;9�\B}u��_5�Kn����뱓r(�yn�b	a��Uz�<�bH\\�~m!������	�6^����F��������"�兪>}'���ށ��#C$
��=�Y���3'Ġ�[VX�8��5��j�|��hx7$l����G�g�ߦCU���=�
���ٚ�� �<�s��x�,����]��!��oR�a��pu*>@���
ac���n�[��k8�=@�o�b�aA�Y��~n����E�hw����^H/u���&�`�EŻ*�A�0WT�l[�M�s~�`�܏m5B���,�_���v�o����/#j��3\����1k
%}�Op��p9���C�4����jn8ĨE���D:o��k��ͥ˶�r	/a�^�����"��H����9�u4^�N��w�& BX���0��wX���gh��#�fo��Ȇ:��Ũ�&��s9�e|�y9�]���C��ɓ�u��B��4����=Y�2��RjP�o��A#A�j��QJ�]�=G�����\�.�o��{���~��w�f(j�J�%l����ј��[tm\�e��������Ak��m:�L��旲W�(�k�}�TTX� �o{XWi�:��~&����I�u�����ɔZX�ԔSu�0a���<�j�̫���wm��"�c����������F��֐� �*FX��\tXZ9�>U�o��9����@f-��C���-z{�Qg��_�$$�t�4{lf���5U6���?<d�񈕸N�$`����ȴx�5�m-1IG��^VD���gg�3a�����1�\�f���!�伜�\���
�Xސ�]Ƕm��m_P�o�K�V��=b��U�fwI�~��m��9pιJ7�|�N�[��ɪ^�dåa����N����'�D��l[�Aw�܏Eu�B��o�#RT(�n}���.���(�q,�@��#2�`��$����v���O���H>b�f$�����h�=�&h�F �N���Y]��r��������1q�� �E��t:�`ߞ'7�ĕ�:<"^7���f�Uj���i8���c�d�u�-N���)�S�-c��v-��:�b��ޓ����Q<�T���c�Y��Ō�ٟ�2�D?,�w^��,�b�S�g
c�Ⱥ/K����g�4N��v���_��jo��{�gM]ϊ�h���1�l>M�N�̔�jV;P!��ԁ������J�SU�e\ 9Nǝ���� �̓�m�j���{�ZId�B+2ݰ"6�"-*��S��b�Ɉ�1�l n\�,L�S��C�x��e.cv�/�ߘ�uZ����ĥ�u�BOT-��"����O�ֈ`��Gy%��0g�9�����ֳ�6~Y��.��B-�gv;�g5i��w��ø]�"����>��w��]֌ԃ�k���q�J�W�"�>I��bܧO��M�d!keo�'���� H�ǭ�<��L"D�������A3��:O�4�O�o:����񊿂�i72�)�N�F3���i�7��ϪD�,#�4�(O u��3<F��|BQP�n��#�>՜C�VX�\e-Uƭ�Z��
�@�Q[�W�w��m�#!zH�-{uW����ټ�ӥ_j���O(��I�p��N��}DoT��V����o˭t9�����yգw���fqo���د�|0�=�a<|G�cS	u_�2՚n;�%h���,@C~'�U���3DɂYTĠ�~F/���Ufޖ��9���Bw.>��AQ)�����_哎�s���i��5[��{ �q�?$�@�^@|WP�o|�zW����1���Z��]��ퟷ���}�{T���1���O
������+Ȓ
�}��L�����%כ�#���
����0�*pr<��א������%'��E�ʀi��4��D���A.��EO�զ0m�bQa�\��xn�(��Y�u
��� �Yux}ׯ�������U�V�{fYmj�d�$��iQ�(��𞎲	���O2jrV�R�_�]�S����Kan�m�Q^���8�v� ����u7��:�s믜լ-���9ȣD]6o�!*�	x|LA(��(�~��� ��\h�g�#��Z��L�:���R�:�h��Eэ{�a#�%�� ��>����I]�K-w�f
*-R�%�v�b)�8�-Ii��6�q�:�ء�|(��W����w,�X+TtyH�j��5������8�Tw�l������
�GN���r�X�2B��/1�  ��3���%�������^o�7�ѯ�3XQ~F:�%W��'{T��V#����Ov�=���ÐN JO^�����N���b�[�v18_���3�<x:��mFͥ�]��2�Y�4�=Y��g=aLg�_������;��o�� [�;xhT ?�l��C/kI���++|�W5ւ��QP�̳Z�M���� S���A�G�ۓz�~��}�P�����*c��j�>��`��W���D��&c9���.n�U����u�*���P��Y 1���w��.S��c���J��kvp�P�K�����xP��/�����xe5�%fML�d���乓r�z:Yx�gcyKO���N�p=XQ���s�:�a���Ԫ�;���,*&Z�0o΋����	˞!s��0�~ ��UA��_�#\G�N������ �0��-�D��mU�m1���d?�O���_�ÚC�c��>q��P�0���,�'�]Ћ�e�
k�h�߱�.�Lȩ�'%K�����0�ͯ�|?�Xਐ_��ڳQ�a��A�tS��X��R r��>dM�Y#֊+l!9ɺ�g�90��X���vAc���h�VQ�Y�溦�o���[�8��1IF�T{.�
~�ԣ<�Rg"�:�f�N�&�����6�W�N��R2c4�4�D�7dCw!l�a��� SU�l>z"��޾^�8����B��pc&�{��c$0[�<�z�!��׹3R�q��P�KG��*EԂFf���8�f�#%p0�Wp�	�'��Z	��z2��Ɲ07"vA�!��=b��t�d"�`��>����".`5��#T@R�4ME�Ic�*��m��m3?x\�i=bJ���}ƿ�]y/`A-7����&���d��۳��_W�ѷ����}`p����V���gr�(�<m�u'*�a�Ĕ�(WN��D����jV0�>�:솽���%��>x�
A�LpuYEp�tx�Tm����KTfj�5
���ϟ��~�9qt�B��rF�*�%ށ��\����:<E�i��$t1�8����;�}��{����&,��%Ķ�������]�ښ#�
%	g.�M�/�W���>�F�l������h>���^\5Y��:�o���prvd"��� �I�V�	_�����O#��ZT�<p�g6�$���AB�=F�B�� ��-��6)���;WH~�տ�Ra��ȱ�Gn���|o��r�37�!��j�ͽ��oLBJ��ų�17���s��wq5VG��}���+�u\��XVYM�}!0���j���E��܊!턹ǧ~a������U����[�ťP0���+�����!�I6�X�ɾ',�;bn~��f>N��Z�� tT�����t�_�!��Fr����;%���([��%�V��+�qfD�9,W�QP6]z�����*����J �����	k�a+��w�5���d4QS�Ϩ�9E�y&��Jq�U�����ĵ�>���!�Nξ+������}��;(ä�i$������1�z`�v��ڈ��C3ǜdU����!�J_;R|N���TŌ�q vS!2�/oR=��z��R{��3��8��'��3���J[��u�+-�mU����6Wu��F�MNC5hy��Wp�?����6�%M�&�t���])������v����5	�g\q��
�)]��K6���w,HW]������s!9����� �
�_1_Lٵ��t�~�a�@>;]���h����PD�'�	����7����@Ø�P*��*&�=�~�9�����E�>��V��y	�є�;�[b5�a�������?ޞf��׿[���q�q �^�!��GL�6��ѐ��a�����K+��	J��R�W �n�z$�)��D���q�T�+Y5����BP(�#��Qu@x�b�.\P��M��%'����0 Ai4�Wh��oq�Q�����P AJΌ	UF��b��s+J<
߲�(���n7c�ҁ�QƩ&�	�����1\�+|g�U^*��y�(������U��Lگ�bU`�>����t
T�����Z����k���$�Gk��zD�79߳�tLU��rծ@iTf<l��.s��B�}��xM�uc#�ې�1;(���.?�����SGPl!y��<,��ݳx������cd�'gu��-7�D�H;���j
x��!��K+B��{H�����z�ӷ,�1q�d������!��)ڟ!/`�TY�	�֌cT`D�$��,��x'eX�~�>�
����K| B@�%�m��'���[Vz��$#y�nYO����Ywɡ������*�	4y��D4�%�����|���T2$ǔ}���%�����+��*�������_#�X��;UdF��D~�J^�~y�T��u��Hss���a�emO�
�c����r2{�y���h E�Cs-4"S�͜��M4��>���ygk<�Ie?mL5\��d�{�/��|�%Τ:����o����>K
f�/�SƫW9\kQ�K�8�o�=[��I����ap�C���
������/�oy��}��),&�!�
��e�vcP�&�lP��g�̡��v�<�;ƃ����!���g��}jW,��,�	�����K�rY�J�rS�"��h��w�hp��ze{S�vV�^!&/�u�Z'� Fql����Y�� �)���	/��e$�t��4��_�ϗF��J-����(FJ@�1f����-���ik_�5A3�Luy��������%�Q<��Qsk�-iF]������y~QOky�'���� �����j,s�acX�wj�N���Ŝ�x4nvpev|�	G��y�8]j��mQ �/ǽg�]�ޱ1Nܶ_%p��W3�~�m��'�_�{}(Y^��|�j�u�&Ǜ�������Ǉ������֘�"
�=c^�	��t�bGo�	!�����jv�?������t���T�1y<���3a�P7�D�af�t�׫��1j�2�i!߹��f*���ӹ��6c#�B�_A�C���y��ή�!+ �	�,	h|���Ȑ(f��(���A<pS�iUU�Y?H۷�:4԰��,��TA@����Ƅ<d�����}x��X����d�7K�+���EH���U D�de�f;΢z��קvl=F��K������jyQw�o�qS?i��)x|��!���\���W����e������{�Af��
@���k��;�P������8+��|����Q_*��e/+���-|�b�H�`X��͌�?��<�%��~I���9ѱ�Ise�Z�?�̖C�[ޅD�cV�֐#Jp�� ��Zf�F�Ȳ!d�^x��;�i~���T#��aݺ�u��=�N�݇���ǿE͹y��6���P<k�-s�Ͽ�d�	4bk#C(�������9�\-�ƨB��@�i0�R #�)��kA���XK�{ˍ�Ջ2�������w ��|<nb4���S�4�mC��������YV�h��M�7b��-���:���'ai�IS�l�(oK>������.�SE�g\fS�Ca�7슍���A^�	1Fm�;E{�N�4�b�j��Ai-wU8i~��j0?{��޲����{]�^�!8�xAfDv�y&�x�E=���ƴjgX �s+����C�st���e�!}�?�4*|f;�6�2���
(2�����eg|P~����C˄�O��fM<����eӷ����r�������\�d�����}�x�h����t�VdN������XMEcgTx�}�5�bM�+���`9P�2΂��)Ѭ?�)���Xd�J����vf�XT�ӯaB�S�Sz2�UsnhA����-:Q�d�c=�&��Gw�lѾ���u,z�}�Ca�µ'x�{#�E�����FT��q}4���� 7��.��M�ف�)c��w�eH���İ	K�o)��3�DX2v�vFե8��q>�k�c�c*�s������v����*�/��v���V�.�$���0�����΁Xn�v�	R}S�P��M����%��B������	��Vk-�ȃ��'%_�?��O��`�b�vfmf��S�ş��C��g*/�¢51�Zjo��p�`",_�<\n{s �x��2��8�8��[����.��w�Ą�2�*�4@�
k�o��,��3`����N�<%t�� މ�.��.�����^ާ1�3f���zW�S�S��|��h�^���d?�* ���?�i{����mƜx��87�#��rrA�.k-��jiOo���Rk$R���a�f.�;���x;Jg4��-�͸�4�Ҡ�'��D�|�\�+6Z=r��5�]ѧ�= ���O�S�Uu6�7�51���q�ZU+M���)���vLL_7f���k��"�Qe�n*(�ɚ�Hf�-���zg\��sB�{�bՉ�)����N�Ґ�P�6�C�$��m2���`�^gO���L�FZ"i$��I�,��o�P;*�i,Kί��dL�[��~z��G��O<�&%����.	��/^h���+zF)B�?�2���2��N橉-*@�>t�<�<���W�,�I���o�K?�k5���*l��*,�Y���oզ�}I��iWϺ�eʛ/BC!Lᛲ�o#t�<�]���(g�ê�3k��?���6�5z0�R�B,�w��W%j�����c�1ySj���J�N��e���`��d,xDU�,�V��~7j��x6E?W�ZȀX�:����>t>mL�5l����o���(XLq�$�U�/=WQ�H�.g�W+��S���	}#����G*�;���,�U&�jXH-V���q�/���3�y�(fe5ӡ�6x��*�HW>�M7	�5=�
"�woIߔ��d�q�A�F�bcQ/!��V�2fk��m3Qd�%C+�e���kx��]�����M@�!p/��"b��Vq��!t���Q�-�E���+/��~s�,��9�E	�7�P�`�#���kW&�޴w^q�Թnt��͑x�u���ơE�瑅ӛ�>�d_ (;0X�c��
+g׻����dv�]
rM@.�k����21����M�*���#����Ɯڝ����o��jCP?�'��Ij3�cβ+�����L�:>�}~����3��J't�fL���@?��}i}��4���Aca Z���X���$�ſ�I��^܇�esIamu�в]qj��I�
e!���'�IwH��
v=����A�6��(��]�����6M�/��?>�
1�Y�7<g��5�{�9p%_սm��y�8P%��M+��#v��;�s���>iE�@��&T��rj��h��׉�����q�(1"i��:�fuW�%���70֒^()R�g "Zx������ꭟ�O(���"ж^qt^g7K+_�o���s�Ԗ�U-hV6��I�u��[�f|2�h�a}�(xŌ�vv��:^�W�<�"4�O��oM':1NÌ�`:��'�.i��H(Ej#��ex�ѿV�����w��=�(m�29����P��ʃ���У�� ��ء���Ю^�cc1��]1!������=Zup�˻�)�Ѫ�yG�m�C���=O2nv���|W���WR�� �k-�G�9�:Ø���D�A�����_�/�ǀrMry�X�n�8��Ƅ��4�&����L���`x���iE2�"j�1���+�UI6�k�i��[t=��>)�?HK�JQ����+���=��.��Ó:��A{+��ul�ul+
�!aZ����hƈ>�[��s?���S�����1�(�)���17�j�A��\���|��~1EW������Bκ1�$�)��dRL8���e]x���a�u���ZV��^��>�%�'����i�F�D�G�w�f��lb4SL�L��CK��|�8/ՇO�	�����-}ʕZ%ұ����f��k	VCm{g=;𣣛���R�N&��Z*�ɾ�~�a<e7����:�8J����=tUJRF�H�G�Ii��n�R�fr�'���(�~�&#8׿�b�\rJ��ХhS�6[V�7�5�ϧZ�$5b����Y )�p{��L\��qs/^X�g���H*+ц��z�[XJ��	~]iVQ98o+Y�/z=���qF%�l��R���I�)� 5�%�,�\`(���-�e�]7V��A�g�}�b�)���з�=~P�/�������pV�g�G?������_6PߢWI/Q�_���t���OZ�����A�ɂ)Sұa�������>n��	s�A�SI��N�"Й-6��S���7�Iכv���ĂPA�*)�w61;X���҄5,fl�Xw�%�PRr]�~������
���/��-S��C�yQ��n�����P�1���B%AA��ҷ������:�r�[f��WVGs�Uq�*׶����l�	�[sƍj_7usH����T����)3�������|F��Z�,D'W?]7��k��a)�IHu>��S� D @~�W����am���5�|n�e�L�Ef�x>���?�<g9����{+Nf�6tu!
#����f_��ч�{�b��-}D��i�ϬNĮ\�w~��M�����g�5�w&����~��!�n�V�*�:���k��Y��n�j~��	v~Wtm�o~\�f簬�A\ߦ� ln���{7q�L���)��Z#����Էzq	D���DV�e��bR9���V1�A?��O���j����,�F�\���np,��)�@v*"�z�U:�y� y�&)ly"�lm����.#�!�oA0Ţ`b�$;$k����
�s=��֐���V ,]R{�/��y�Ԏ������|�1��+єdT��g�,����,�_���)u����R����tf3Ab8���Y��t?qs
L��̿]�/��]&��[:c<��؞�(4G���)R�{V�g���ȸhp���YG=_H�ɐ`T�!�P:N��K"�P*�A�\5P(㿺n�e6�N	G!h��_"�6���H�y�O(k��dJs�贌���^�9_ʪ{4�*W˄�;�x&uj�v}�����b�-T�q�@t�݄�zq��(2��j|��`/� �t$XR6���w��K���5�ɽ�����e��i���X��IN����=N���Ǵ�L�
�����u��b��Cl�v`��$�}k��&��|M{5T��B	8��eὧ��%q���y����� I�� ��,lkV4��͊m���G�ϖ
,�q;*�E"W��Kk��o��|� (NYw�rC�;�s���z�_
�O�A�Q��ʮޮ���lh�\½h�v��2]k�X5�����Ged��b��:�-�=/:rg����$c\,ɲs8��$틎])�.Cjv�pa2�;��� ��.���p�t�z�
��9���#V`?&�f7�N�y�)�=���hjN�E�WF��u3@�;/��Hf����`S_5� N�S��DL=��02YE�I�N��8�C���8����9��������{ZG�U��tj�*�b����e����T*㊚_/�.Y���43��c�QKT .� H]m?�� O����ag���(�S#��Q�I$D�6}:z]*Y�E[�S���v���aZ����ZG� ���5~Lv*Q��Ӏ7��������"6���?��n�\�T����Z���3��%�B	3��]�5��8ɩ{���a�<*z#f"�� �^@�H�������U�~�b8+p���U!Gf�D-Y1�<d���_���!����4�ԁ��PX��ZxC�_'��{^�Lq�R��@h��me����9�.J��@�l���p1��`0�rS_�yؚ��	\:���O Z�aR�����s��'��	Ä�vxʊZ0�����{w&{̯�{Zu(Mm��v�ܞ	����� G�סIx�}߃��NF;Nr��[�ymԏ�%�5Q�蝶i��_�{a��6��^��T5�`˚��܇{�O�x7�
�����a� ��jb8ci�;t������o��k��1â�-��	�+�ӵ��8���i<F���$�;�Օx�x�,-o��
fޅ��diT�$��_���8��Q�N�^X=H�T�aO������g4-dk�g���,4n�-��!���ܸ�!�|�9�-�/WG���G�{T�v��?��RZ|��_��-"C���:�>~ʺҖ^�΄��$~)/� /�J~��S�Hg㭺�M�;�Ѧ�o���#���%h�6 �?o�s�?啰fq�ތ�Y4*���ub�%�#Έqyx�,_��[wX�Hf�-�aPuTO���rɌVM'L�`hH�g�|[�,�ӟO�Λ,zĿ2MY���Z�v�NH �Q�GW�E���-�t���YÃ�-��췁�_�$�qD���<�Uqo!�9��%`9d(��Bl6R]o�W��G�'��t�U�a
�b���(�2���o|�-�5���-%��ZR�Rs�U�A�LFdn�
���_��f�d���Q�;2zF	�/[��A�]��[���t7\��F�!�+��y�7T*�|h�p*�	@�o�����/�Ƙ�	v�wr�MSaaT(ݶlFn�I�-Z�5Cy zBı�����YF˾o�=h��V�l94\P�`9̲��kB���4�������` 5z8_{�>LnYtC������v|vd��ޝ�����<��pBW�'i��`-Ќ����y�����J�Yc(��}����_˨�Z��q�>J�[/�@�%��	l��o���x;�͑�.ρs�$��7-�H�XP��8KC�Y�[�fM[�VOȎ�����}�V��w-D�%���(~Y�6�����c�J)D{��c�a�� ]�����5��Ǣ���;���k�m��v�m�l�fH�g�dO��(U��7�I�}t�Y[<��q���"�T*������Px�cC'�n�%�ǀ�T
��v�i\vC���ľ��/��!n���v��{��Ǉl[K^BQ�#��a��z�=��h9h�Qd����#����E3�d֊{���P�B~��F�I�@���_Mp2�ɔa�"e{�.
B���"P2�Xr���3��6r��x�'����]�.�\h��j�O}�>��vZ�^w�*�i�a�4i�-�ٙP�^+� ��j�o�̬�.]"�@�Ag���A�\��!�1�m�-*��V���{�\8�>=_e.ɶ|�FmzL��\�I���d#*��
��?�fߐS�w,! zbJ�L�J���V� �+���//����ȱ��lAE,�'9�r���k8��3ȇ�z��J�U��{�MG�x���F����_dY�1A���e��q,�Ԯ{;JɆ�~�};����}���#���.s�l&��w�!�q��65��<b���u�~L�ԏ��K����Ik���/����z��г+Ҟܮq�|���#��Ձ�f�,�+�%L�,�w�l���r�[��'!@��u�{+X�%e�A�aL��	ozY��;=�W��ۑ�x�\t6Ύ��*���8̓�}K��݆�~�,�J�%�C���g� �
��O����M�k��/�b1��*�3�ӏog���i7�E%��$����%��8t0Ƴ�Nw��i��y��NK�f7�#G�=�vR`�cX�t�1���S��6�h�udƜ�`�. L�;�􈯔q�V� Ҕ�j܍/�+<�q;���s����:�a��ǅ�f��2�8���9�әy��*��j|L��鉾%�*hF^��-���Wס��_��`�W�)-K�l;���.�hW�5A��;��H�`d��D��)�Y�1��f�����_�`�A��(���v�q�q ��4,��9bXb��{ހ4B�$�4���c)=�M��!�P�p8i�H��4N�3	�e+:P��[$�s*9�[ҫ�V�^!��f�{!����F���M�!�q��H�"ːucL-����HGo��0 �P�\29��ZH�óq#�q�EaR�,�+��V��+'MQ�*�����j�kc�Q+��8o\��Kj߽�r��0��Ud�~�F��we\�^u'��٢�Ci��o$�L�P��+uq�A��+
��q�;y��ԃ�\g��sD#G��#��"�f���;Bne���ѐ����	��R

�DP��o;�����5b��Wf��	�����q'jh�[M���﹪0X��.+W���=q(�T�`��+6��/�b��kJ��_�� ��E�g/�{qd���{�aI\��	'��S��ZH�)�:�!ɥ� ��[�  �fR�-kV��\J҄�q��*:�s	O�%ф����C�%EϷ�#!��7/��ɷ
�Éf}^3e��j�9H	�  �8����	~%�a:[�I���N�*|!��đX���9�7����g��瓜���M���?��0�f�ol��=�Sι�Ds�XWs�Ƥ�"���6ows�D�w���j�R)�`�w����UJ�k��>x�X~q)��o.yV���і!	<�	-�&�`���,] 3��t�ʿ��^�y�ꏌ�\4a�����Z7L�*430$@tO�Z��:3}�h%�i����O�)�/4%�NO��$sqK��|42�\�S�v�ȵ��D	�#D�>��A�6:�����ֿ��a���~�j<p��)��7z��^����ʌ\�����s���+U�{�m��\�~�F��0�gVo;�9���BI������|
���E.w�[\��PB��ꘄ��e���Vԥ�=:���0= �U��2�9�׺��0ӡ�ֹ�B��B{Ū��rubD��F��1ȋJoU�i6����gF3@���ݘ���D�w�a{����T$��p��؀"��?�U���x|�W�e������c���o�	ABW(���qa�l�����9)�[�yj�th���e������yZ_PH��\ODD�m��=�G��0 �<��G�������g��(O��|؏�	�]9����3�mRw�8T�)��S����g�hZ_��8�5��k���RV����YBJfP�]��%�٠<��͡l���Ւ�{`��n�����E�+C	_�H0�O�uYQ%aA���{_��U���
2��|��*��k���P�c^����]@�Je��<lH��2�̝O@_�o��\���D�n��E��c೮�L�a�r~L�B(Xa^|�"s��tzZmܰ &�G#�������,�:"ݤF�D������Կ�����;�p6�Z�ț.H�:8�t
�w)^�@}r�3���QY�/	�����ڍ	��Q;��o^G���!Qˀ�`�;$����6b�Q(X�i��ͺZ�	yS2mZm��=Pa�rעɪ��ݼ�����OB�r��6�>�A	���������>�w��ܞ�υ/<�������%R�c|"� �@� @��Jpj<*!ϟ`;b,|�x��횔�uOcK���v�@|~c~������iBA;�QT~넍���]0wU�߁�8����!k{U ^}���\��w�Z�6���C"�zy����� �7m���M���r~"$��O�T%�OjM��	
��W�=����&:d��2�I��L�/R�:�9<�L�����?B�����%�C�:���df�0��Nګ{������h��(}(fZ�<
=�"-�ƿX���.h�e*���;x)�l���C����r�ψ��ُ����t7Hﶳo�bɁ`�)�%߇_~�IІ7��;k�g�j����ԚP?R/1M4��	�G~�.�W���e��e
&��n�h�Ȣ�L�\¯��K�C��a�	�3>^Cz6�8����c�=׼�.�|f-o��{��4��@�/}�`�Wᒥ.��C�1�W�qʞ�)�`���LL�fZ��!���U����md�ٚ�.��U����G�U�b�K�3w�wO��s}״0J�q�#�'F��_i��[�Ghw5�d/��iuDJP���h<n>'�Hju�EZ���_�;�zKs�4R��-��]8pT��ul�.B��4�E�x�U6r���������7R�O���jà(T(G4��q��a�OɃo�m�;\��ҢݾRWk�K��4K�s1���LY�������z��|kA�}WҮ��Ɩ[��"50��ͤ8;S($�M ��(��Q
`�!߁�*/�������K����'�4�Z|G>�7��Ď�AQ�yk�����O�Qy�2�b	P��4Y��QW/m��V !dɗ)�S��X4�����p�8�4W�d��Aٍ�Nia��E����7��=k��|D�� ��R���Tq��wi�)ݘ���{$����3��� b��|:f��۾m�y��w�y��[���{�LIo"STܽX���jʂê�z�.D��ʜe���o�,^�D��c`�vg��:/��~�G~�v����Sl�^ʻ��YQ��H/�ֺ��@�
إ��Ӭ��t��x��ؙt��g�̷^�tv�%����Z�T���[N�$s��G����oF2�Zz�+�%T��j���]B 2�l�^Bu�ޭ������jhJ�����ؽN���q���O]��ߜ�'�c�m�L���H�33hV�-d
҉n��7|da[P�֐"��JzL�Z�z)ͼz��i�t#'����t�.���o(Ò,�}wN��i^��V���`�-���M� ���9>aG�A���GBX��3V�\�]����:�R8��'�.�YS&�Tz��]η������5���#�h(�Z���Y�<zk�k�-��'ғ.�zY�x붎*�y�+�:�]����T�Vt5=N�u���{�(��T���2\�r9�<��>p��݂��gX�Z��y�&(�Ȕ
C{��4D`Do���a�c��;s$�eꅗ����<H�5�����ޑ���S
.GO�}���֨	׋�LP�j������1��|����~�EIV�z/��!=��a�i=� �C(���[P��r$���J2��3@��+�'�k�� Gͣ<ow�n�o���դ:��x������FxyZ�W��'X��C凜�l�og��uc�fS:���(� �%�!5}��Mh�ʡ�.�*��Ϟ:�sl��ښ
�&3�O*N��b����z������!���sUi�M�A��K�|�!x:��ga����a��.	V=_Z�^&.H��F}��mim�q?��9i�a1���|$����Է��?�iJ���J�r�e!PJ�ؕ�uRN��(�#,�޿��a�Y�v�S��!C��\J>V�����gy�ہC+���/$j0����z�2γ�4�V�E�@Kx�݉���������oXb8옠�~���9&i�_i,l=U\�f���A	��������c�A�?��ݣ��1,S�S
tI����]�|�w^���`���v°�=��O=.�.��ʹ�������Ж`ڵ�F�m�x|=g��q(�`�yiz�._TD�n���c�1u�ި=���[�T"JX��!#�Sէ''�v[n���Il=���SÝ�5&��n�h�bN�Ւ��K�j=��&�k$=My�jj��"<2���:��n̸��-�h��&�����۸��N���e�˶��7��I>�q����@:�ۄx��,}�ç��٦m���뉃0ڬ+V"�s?{6Gށ 0<�&5D����7^�"��`7�h%%���z}�_�R(K�`Xb�$���Dt�G���?��v��a�5��ɶ���Fk��`��B031�?���?�N����f��,�<�xVn�R+��,W���x$�͐��u�@E�ӌÈa/��
 g�ɦԇO0Se٢�.s��q�m����[��|g{�����gXIr��0N&1q��d��Q��w[�#�%Y 2�EG$�i:�Җ��S�_��}X�΍�i@n5X ����-3��끥5�bRʙ���̦ ���XU	��*BR��d<�ǋ˦RK�>Q�Zn�^U���%��@GḄa&W�>af���]ҐO-T��Fx}U�3��\j1��v�fI�al�pa��ef�N���"������)�e�8�!hJ��i�Na��-����'M�cX���r���ڇ�ψ�PYi$̛���"�7����I�J,���
'K|�Dɓ�B&w�Oܯ6�ǨBl��m�tdn�*Ȃ�K7�#��Lo���&��r(��N;O��6�0�D�kՌ3_e�����)��9e��ꤟ��� �sKxdU���R�eƏ���D��bf��a,�� T﮸��&Bcy��>��w�O<�@� ��e ��j��.�bf]�h�Ə��c �g���~@�����o�4G2�p�A�6�pae���B.a�ѷl�{�|�-�du��g�$1+�مx�b׾[��oR��/��� �7'2����9gOY�c��*�`x�ky'Ia�A���=��0Ɣ�
ur|��.cиPQ��]5�yE���C�ku3J������!$�7��c��'�+����}ȆS<��aW N.�񲄉�׬��:����V��0,�J;�W�L��H?�A�d9��	����okMH��ID��A���kֈ-sy��7�P���GE{����0Sy�����%,Q���zT���p�h��qtDj���Dh�,��F�#7��r&�ԉy7X��X���I�ߵ+�P��-w�X���	[�X��w/�'���$�E�j�5�`�!�f�*��/y���$ɉ�4$ Bk&\�T_7�*I�-�3[���%EV�:˙��l��2��=�д	Dy�Q��>{��N�ôV������J��[Q"���Csc(�I�����$�T�� ���t��|�;�,�_�9�o��7�c���n�G0lI2��YƤ��	zdF����`N�z>�������L�o䌁x,Q!ڠj���"��㡙o)LV�1�ׄ�_�)����A�?��od��0���\�K�D�M�-q%��?��49!FZ�6�ąê �)A�"e�[�Se[cƩ�h�rT� S��c���uka��2ǬY�w{(d��<�@Y4|yO>Q!"{�ܔ�f�1�*�x�P��2A]����䩸��7z���O����ys���\D�j�pTr̹DQ�Hι���cQ�FA]�?Ɂ.��r�a�8��w
��J� �����a�Q�n�J疅m����:�z��5����:w��Um<Z�)n��~��8m��ۛ���c���z���ܭ���5N�C8v:��v� �@�}>P}��"���&1�t�I��b�V�9r��a*V�����U�ɍn��ݤ������l�����a{"���17�%u+�P1�a�x<,�贑3�2�%K˱�7E�O�.��=	�+.:��f3�s�~
Ч%1FLY��2-�i}<�2�O��n�h��j��d�=S�c��:s<������� ��L0��޳��>{������K�m�Ǌ6A�o�!Xu{�G�\C!m��}�O���I�%<�|Y���/R���\g �״ݼ{�T��O��k��-�D��0D�hf���W�A�W'�����(3�@͐�{�sn�#�w��H�=�)|��5�1�!���ew.����������QR����Ɣ�t	�Ogp� ��6��'���e���2p�sT <*8��|)��4��ze�H>{�L����FF�<;�ž]�<����n�x�����"S?O��Vhn��I�й=QY&�$�f-�+r�Xc�M(�ݔ$���G��$�3�a��Z��r�G\��uN��/��K�s �sEG=!X4�]��}]/7C�e��I�ܕ
_�x��j�OgO1�WX��V��Y� Ԧ@Z��l��v}x��:�2O	�Z:��j}*��S/�ek�_�T�qJ���x�O�T�3��6���"��T�ҕ��B���*�H�{lRc����Y$b9q�Y,*9��סj��{<���5́!�K��r*��9�g�߲�,_�S�a�w�Id�O�ؼK�����8�@預*�8mW�"���U�����|�3�b�B뎹 �mf4,�<@M&?p�Ql�5��߹7@���e�pd.;��7�]fi���,U$ݔ1(����uBR�Ĕ�z��guh}D���Bx����6�1)������6g>�H�X P��xMul����S��
4Ey��u��.�K�����o7~-lTt !�l���|4�1�$�|T�I͋�B��Yf�k��@�o{\Jr/ y~_�wـ�C�Y�6�Gש$Õ6�����&@8h�+Y��j��*����oK2�qI�8}你MM�W���]e& ���7���=����\��y#j΍Ш� 
4H����eBn���4�{f��4�c����/Z�N�3���X�DF T�,�SVgN)K��Qj}���8�Q��!L�F+�*�6��>�F�(���d5�7q�7� ��=��
u��U�Q����o��
��m��Z����n5��=�B�\���I9�P�N�i�N��݅7�O�P�N%��8s�9�2G�H�c�T~�4�'�խ���H�Oc��?�Bh�=�d��-�*[��;�b��D�$�6*�>��z��g�c^!�Z�d��C|�ы��r�er��M�IH�dbr�uvϓt't��0�AuT�Sּ�\q��������ɣ<������0�;.����oQ�?!��񇗟p[�N$��/N}Sm�{CS��!G'��9�u�z"x=�y�f��g�0��aS^��n��Y$#7�y��|��l⣧۰�tE=T�Z��^珷C�f`��������l쁔���Q�҈�ٴt�z�M��e�fla�BG���:�	,\W�A6pZ���	>0Wfo�#���NP޾ˠ&�g���ds�5z��We�
�����g{i=�����[����g&&��ho)��>��9i�ٻN+5�|Tr�;�TZ'$����"��ȢI������)�i����\��?�czSE!dj��%c(��;�*e9��{Rk���Mgf���Yْ��E�4�����w�mvk�w:�쐞lI�ZN%fF��IQ����6�� �I������%6��}Ynz�ݳ�+JP�8\���h$�x~\/���(-5Mm��X�`�B0�Z����z�C�d{7ڈ{;$�O�@NVikwN����)�^s0md\�|���7��,1�l������.䖮����h'/��ϩ����aP���.
Y`e�1�g���"�r)C����*�_$ 'S�KF�r������۱\��G�A�"�ؽ�l���H}-9������K)ͦը�2�"�3ߣ��.��wz���@�P}�`�|��W@��<,yP���-��Ր��2�wʽ?�5G��Ğ�q��9�d����1Ȧ�8�L���H�⑬���ʛ�z?�m�G�!umƐ�ةW#G~0|�a���Nʵ�m�� \����+r̹](�_అ����vl�i�>GG��n�%[��A뽎nZ>6spf]>�D��R��5��D${�K�����Xt�V�Ҫ}�vF＠Ed&��H�{�:֓KSoʲ��!P5>N�a#|���𜿗�	}����˷y MZj<����0"�J�͇�;j�ϣ�u +Ļ�C8h�'ͅ�H�6�����W{M+;䭮4e�$�����s�Y�P�kW;�A�?��1��7Ҍ����ۓϛ����}1Y\��<w�3/O�ڂ3t��:���|19����4#�`+a����I�˾vJm�Wm2�vVY��Y�����b�)J� �祴�D:�k���9�`,kH=�&g��֗��N���_��,�*����-�,����\�ƁB����Um-W3���FL��3n̡	W�DWOG�c2����Bz�Z��C�n1�_+e�(�77g+�|�N�Ew�BZ�|�/��kq��e����L���Av@�(�N�eG
�g�P(����ƓtJ9@�);�w�g+#��á)ޗ��Ǫ�l���I�>����Q�#5KB5q�>!f�i�n���ώN�t���Jhݺ�ԩ:$��aP�a*��R�c�}or�>�-K��n��_�*0��J�!��`�JIȥԼ�;���B��DȦj��}Ɓ��$)h���Ґ&w��"`]���%� ���N [	�v��xM���ԗ�jӳ��غ/��Z���s2�Xd������8�L/a8������?�n�����c;�׎5�UQw��T�4����.�C!���| gK�;��U2�9�����rW��kY�w�f�Y��\dUr���ؼ	�Ɩ�I����w���t^��)|�����E�K��W����'>�B��ё���-$�}?C̛�t��G���Y�t� ��d�>U>�w;=z�>f% ������˗���W��{&n��=7Yp�Eu�ڌ.g�7H�(�3y��1��B3Jtv��*wgݸXl%E����&�C�nع���Fu����@��vʠdu"F�a��d<�_��QXy?�B�U��65�qֽ0=�$�ؠT�z�����C����<�詻⎃�M�̦S���t�3����]TNt��{�r����
mvЃ~C�a�=�ˢ���F��|�����H:�b�7K���!���b���|�3�d]f��F��7.����e2D�dAX���+�s�SRN�,��;�+8z�W&o����ݗ��ø�Ǚ��L(}j��2�B�	ɀ��3�%h������H��$<�����!�N/hjEmU-%��MB���hR>K�?@���x����������.ޅқ�Mk��+�l��C�����D!�.�?��1�/��2<~2-��eK�>�/n�x�'��"�p��yn�,��=�-1w� ��&ɑK����;��T�Ю����Z��2�k����'��Ol��.ġ)H�X�]ba��U�:��i�l�m�����kK�~��W�^F�������*��ߪ#�І�D/zw�6�@������ТM�|��&�G�w�nޠ��Y����r�@�v�W��T)�ϯqC?��C@F���_~�!?�\sz9%ʷRH�R.bb�#�Iz���yH-�9G�^D��{�}��H�-u��+�i�F#q.-ߏ��	.ќ��5R��B�o�B�u9�����A=��*�a|�L1�f����W)�M������6_Ŭ9�����Qõ�n*o�B��c��޴�xX}��f��-[���ʾo� ���	ٚ�Aխ�t�5��b]_��i����%/�|m/ܠmZ���q��ς��iKM��0n�<?��D�5˷ ���A�k���Q��.|`�Ǯ�&��S.�;�VP��i(�* �E��j������Hx�ځE_C���A�)E'q8��	�2���������hH��N��d����*<�4����D¡2g
�2q��׹I w�������qDb��zU��\4��$]r�fRoI��\o��jԬ��>��:�X;s-5���[;�m�B�M����r,�A���T��㘛�o��t�����9/[�P�|�y��TNB����P�c*y��uCR�-��}Ԧ�D,-�c���o�x9�2��j?X�#�n.A�6�8,��Ń�Ź�p�\tL����M����y8�Q�}L���Y}�
m�B��t(0�e�^80j��bMiNd"��W����)����F7~%��Lc�D=S:�vb��*o�b0L�D�ї��M3�L~{��,\H�iU��s�n��L.�Q��p]G����][ﲬ���VC�V,��1��\��i%S$'��1-Y��<h��G<�ĝ8��?S��^��P��'3Ie���M���3��8����U�� r�d�T�$�-��1��46��, �%W%��]�d�M4@,9����Ր�kTX��GSg��k�2w�ĺ��l%�Xg!q9=�\𴨐�-��_�0k�����^��o��8�מJf^9b�10��|�����{*���Vg���N$r� "�?�h���lM9K�E�9�b�X�����&�<nE3���.�J�Y���6Y��i�o�,���6ƣ]��I�y��'^��R�W	^#����EO�k4C��]�V���5ϱb ���u��+�R:���j����cng/"��#�Ƈ��e�"��HV�@��/���ZHo�6�R\���Ȣ��;����	����G:���G�܌ы�d� V������d-|�&f�͓K:H/�ɰL� ��gG{f����-���~�ψ����'&�X�]i�5.����W'c91y��~�(3�՝�P��K�M���+�\O����d?p����a��l̈O�\P9)����g�e�({���@2���ƾ��RM�r7ɿ#�4&�Et�yK�� �����*'���&��!-K����~�^+�Q!hĕvQ��NO���� ��奈����"K0�?��Z!W?�̓fK�2@�-$�^��5#ԦAߺ�r�Jf�#� NHZVN�sB$�F�Ct�n�B��8,'��W���4�Ŧ�l�f�=h��T٤LU�%jܐU<��(�"Qh��b
s�T (,:!���cU>)�kw�n�
,����I�;>@؄E��D!����\�� ��^��l����K{:�f-���)�7:pX=uY6�kc�I�D$Mwh�ˌM\1�K�kεj�V�_�By~sq~�cx�J�u�_��N�L�w�WK eW��2���n����g[�{�B/��t�uM	���q�/�%[v-�}�jGZ3uD�a`��Y�v�y��7SL�D��q�$��6������g�� C�� "��\������ȷ@��s+��9#��~���Lt���!#K]� ��d}Q7թ�0����ۛ��W��;^ӹ_�I4V}�:�W���X�i-�ݤ	�eM��J�ܬmp��R��!�@X�`B��q��U�Eo�����	��!��	��n6�M�>5�)��a�a�@�n���(���>��A�1'}l�s�f�K��� �6�ϑ�ě��i��&��d_٭���J��Ѩ�UI ��,;S@�yچ�X�s�]|�/裡�A`��,vA6ddg�=:��t���;т�!Z��Cɥ�x��ȅ0��4� z6#��X�k~"wȠ�W����S��_o.� $��C�����C�}�[�/�/úʷ��
��k2f�2`$�b���"I��4X>��߀NS�F;��O}�H&�̘u�z"e��w���Ɏ����� ���f�_��Mv�sk������v����i���?�Mw�[g�W���{/Y� �/����0����JhI��}+X��f�[�Q��œ�G��Z���-;̙)�J*�T(��x��u���)PE���a(d?rD|hEx(��v�j-Eĵ;����8f\�o�y`N��1��T�'Xz~:%��C�sg����xe�z�BA��o@�<���t�Q��?h$��5��`x���TҞ5�l�����(_��){��m�$�I���ki�� 6�����I4v���eW��D��>E�G��$(�0?��.&�p�&Q��H��	��n�]���64<�_�?�Bb-%��|{3�;���߭��[�B��� N��Z@���3���d�e˄Vf��p�O�m[hX ��m	Ա�T��d|�U��軠;AgD��L�l,��X�Ki騤+s�o�8㓲��Pj�g�%������~~�v����ro?tC�>�l���G�ج��i��;�ǩ�9� ���  52.6�����~�!8 -�D_�̾��+��D�8�E� έ�e�P�1�����f>B�q�������(E2hqv�.;=+�,Ќv�/s[����t)��
���!:^����J. v71q"p���� ���`%HO�R'��a�~F(۝���֊4-w�ᜟh#��&��y�F����pai�����
�5^�)����)�����`��uG_ ��ɧ�C�j�l����7�4Y[��]?Y�c��V�\Lx����6-+��f��obr�������v�raF�6�)��,"��Ό��(�et�wDXɰ3�O3����ra�Zd�#�� ���U=��!hE��n���gY+ě��-�X7�&m˰0VO�}��:E���N�~O�N���W�&�/H�i�֩&\	g��5|,�(�L�Ie]���/��HcR�f��
�U����=�z�`U��I�@�R�cI<��p�T!��j��"����#&f�Ш[K5�u�A���`i?ɼ%\;��ÝB��(i0�n�F�:	W}/�z��I����|�P���Ÿ��AKx��و���	ZL�'f,��RW���i� �!7>����`�A�����rG�����D�k��"�Y��B��9;́3%��6f�7ȑͭ���^�ak@X�x����8l�?��
>T r��� �.�S��K߫��)�dŧd0�|?�\K��[�H��WL�O
W0�r�j5�����1}�N�o�-$���2a�c&d�/2d�(�RoxH�r�h����$�_�S�pm>�����VB�Y��`B���!�@�'�cdج7��[�#s��]�t���� ���>͵��C_b���R�bm�_�� ."Hw\���Z
{���&�:�cvrT9���9}H�<Z�)lYU�!*�Ö���/�g��o�ɿ��"�<x(Z�NaQ�i�P��Y�W��v �Z�>0
�!>��:�%��z�d�O�&��T>,�]�:� l�ޑRf���_D�;���E�,��@&��(2�
��b��cGG/�]�g��'��<u��ޣ��R�P�j'Y���Z�܊��Qh{|�u��)nJ!�P�����t&��U�]'#|`Z�o�Le!�5�EV�5�r7>�]�Ӑk��o������[��DV��FQ�]Ϸc]��4Q+)K{$��{gj�������&Vzn�kCP�nx.��B4�c�T
R�ǥ�ǲiz�L,Z��ݳ'�~�Ơ��z��\�+�������{Q�YE.Q�W=�����U��ہ�J�7�SuS���i(r�+��$K��[#.'B]I�����=�j� Z�3~d"҂�m�Mm���X���h��󱬼���x֙ ����9�����AE�y��Vò������bz����X�7�V�yc�����8�
a�!�d7_6�����5��/�0���}9~������ =����X+���!7m��+��b����1$�^v |��f���eheH�����n+�Xԕ���W67Q�P�:(r�tѵ����F����]��w�B2�޳RCr$�e�9�~&�?���d���:@P��a����'<���P+��ٍ���j�!ꚍ����� �W�ߍ��;�jШiK�Oerє� gN~��Lrhxo�v��������k��q�x��ĉO�ԃ"��M�����&T�K�'y4B�2Y�m&���=����֙znS�������>&w}�b�����wիB���~I~���~BHg��s���n��6���aj��VL6�h���PD.�db�.��YQ� ��C���rң(�-Im6�`�� ���dAO-H�؛ڒU�7ml�C�Gk����ʛ-���z��d �w�x;O�9����U�y�N���^��M�_Ť��ǚέ4�lHDT�1`D�Q���Qb��n�v���kt������(��<Дr�4Y��!u-��\4��A��l5��虐�S*e(�<1v����������鉼�#�QY���'��9.Pw#�qZ-�Ԏ�d�� Ҏ_� [���3�kJ����t���@NK��Y3M���8R��03dcy����}�W��['�){6��k^���z+��׍(�;Gj̀�ӑ�?��o�am�9�}�@��
�J_�)��f��qf�Ş<#4�X�O�Ӷ	bLt�P���*v+�3߆�5�H4LVG����6x:\���~"~M�\�'���[�yIDQ��"�@�c<9�2$�LA����ӓ��W�#,@����4��"c�Y�B	��䠭���l�x�^���B[�p��VnH���&��hA<a��ƹi�9F5E�g�N��̎�x���$q�s����1�i�}:�脤4��u
GL��9��z_��x��t$]�6�F��ǡ],_"N���?�*���7�����@Rz�E��.���%��d�3UK�&��hb~�r4F�R��%�t��S
䢄�63�����vg�D���L#fX�x(�'"qw��&���
���Z��?`�(A@l�m�S}CS�k&E�ْ4	U������}��HSd��]���Z _5�ţ1E����`S<-#AzV�t	�����k����"ZMZ���w*�֫�{�
���#���d��)�7��ө������#
ş�&�Mw�L�%;䧳03vMd~N�w�r���x匄V�(�� ᯨ�+�Zsc؞���������)�dM^ď�ˏ�^�S�]�w��X�>:��sj�$oh�z���*5�7�P6���Q@����c��5�90�Y/�
��}�m��n��W����"�w �$�>~�>8��w��Y�y����t�Pt�q�4 -���:�s�%#��SvG`��Ӫ+�"l-BD� �۶�KZY��#wl�g�Z�;a�иt�P�?��|��zv{�%�{l��p}K�x���O�/���ٷ-t'�51�Hq��X��;���$�3)
�ڽ������	PD�&���**�������������C�gg�o0aED�N;³�qM�ӽJٲz�.ȃ���i��[GW^����K&+o7+Rؾ���N��k�������#��㤜m��5wP�\�'ÂL�ZǸ2Sd�_V(5A������I�c�4n-��}��{r�7(Q�X���Y�5�;c�qO�ں�P3=���@�]��Ȟ�=v��T�vu���>\�-�S/[�@Z�o��!���J��_��y�E�qF+���)i��7���}@b��	�
���N��6ʧ M���i�nW�Ǫk�UsY��	�������v���>��>;�>r	䴞���q��G��4�u�g��/u�~����(�m�K/���ӆ�B�����p�Y���Í���x��`,����:wdI	}�;g�Of�Д��+0��M)/�U��p����L�'l��ܭ���Z�H�(�B���sު�Q�z$����B���8����֫��(�fC@"�;7�z풩�D�"ԑJ���|&1�w�$W�m��T�H��wkV�ԋ�q�L�Í�pe(~#��+y�3�1-��8Ƌ�ѧ9jn~��%�:Ҫj���X��c���>�\������Qɘ��G\ZԤ˔wԎ��ޙٔ��#���n�N�ȑ��a���&���ƏG+-�L�Ju�V����x�n�>��S��B?h�����������>u�ܘ#��GdM���-}�U�iO�ٕ�=�V������o!O�`z�S��).�@�cG>p���M1<K�-t83�
ə��"����w��]�ns�@u����5��<�<����N�����*x��-�j��r�à+ljm���J�Cs�C[��R�+�'�H�'�A����;H��
�; �m����`�/BB���hzh�&�	����f͊��ND'��3{�G�:�9Ԡ'	)���YB&Y���R���&E�q�l��<�r,L)"��,'���(���Np����,(�#�cs�b�ၩLH+Eݛ��{A:��ZlW@�MA�a^�T�lw'�_���]�ְG�y-���PC���1ZJ�8�=A���2��9�H�����ȕ5Bb ���v�MBꌩ���t��Yi,Rm��Z�CӪ���38�δ���P"���I�������!f�cܵ��?bg�N���;z9*��fV���q�<�ڧ�ȷ��C�ywӐg�'�������A)���[��P�Vk�̩�_��u"S�N߹{���4��&� 6�1�n��W�'�x t�g�,���g��2v{~��98�[N&bض�xiԸ��K�";��;�-�8��=1�='5l�'�о�D��S{0�I3�`*����I�����i���#���a���K����2v��p⨶8�%w�zJr�`��2�%����)&�{��;��H��`�b���r,!�0>�H���4TjI>I�#L�]�c��*#kv�#�-�t�:�閹�{H��m�B��(ܔ�ǩ����5ä��7s� ������hބi��d�����ԃC@>�<�ɲ�.��8�SVqnY��*�t�7�Y�A� �6΢����_^X&:E��Y	4�����/ؤ&��Z8�SO������_`����Z3�Oˋ|�ss�ip)��[kj�_�ڡ��Pk�]�J�@��!$қ��8V~L�99�=�5�}R��J%:����1o.�{�	�����Q9�!FA���Þ_L�6P��Z�.Os=����~<Jn~�W1�-]��eW~��F'b��<.���˹��(�R�!�zt��W+D弁:���x����mQ�1�]��癠#�	卑��Ч:p��@��Xn��,�m�z�|�}hy.1gId�=ԣ��J]'��U��+�ԇa��{��~�R�d�4ҷ�A�y��A#���B���E�6�cnɚ�A��zP	2�� Hh���3U���ܵ4��agш
��Ḱ�o��o�l�b�V�e�z0���)<��Od>l*�L���S䵣�z#��	�'�(����}L"� H�,!���u{^�d�̀A�gC3�=�r�aÙR�ߺ]@Ia�k��"���?h跰X⿂�v�)�t.?���<�()���D
&<l��*�0�V`p���qb#���A�0gZ�T���*��o�%��Y��/�n^m���z*L��=6<�4����<C�E��e���5v�dڕ�X@7�O��g��@sv�`�+*#�G�EPO�E�<h��Sc������&Y��v�,��J�������\����m���2%�c��Zȶ���Z�r덒�~jKPH�hbș�'�i���t�?��?E9���Dj�����z֮�V���h���,K����N	!����pF��~�;:�N�����H�D)��9t�S��QF)�Moզ��"�y'�_�[�%^��	�˹��K����v�L(�e�[���n�d`]��Xr^|<��.ξS�U�.r�Q���ʋ�:��.*��[���ԝ���q>c�(y�yp���0X��M�T�ȑ�d��(}�ǡ�D����xIk�*/�ū�����?��zT$8�t�Xn-�o�Ӑ����j�M�����هr�|��C���)�[f�&�$@�V�T X)U�t`Jj$�����Uި��N�]0G!����R �`���c�5Z�#��ޥ�D��Ȁ �`�}�T����z�sX��b�|��N6iGav��KR�MA���ӯ].��͜q�W��V�o��D'ZC�E��yt���tj�e� ��-�� �]P�f3>\�(����Dɾ�A̘���U/,!l��䥀3���JC���{�>;�m�l0�C�ϛz��B��Ao�z-+f�V�b''��-u/�/��˱1����ՁH(ZB�.H�A�T��(.�B��҃��6s�:ԆޢHv X^�,�fy��.��G���p����@qqP���.Uh���̑���}�4.���B۬����Ȥ�Nf9����^�U��l�ִ���7[{��t<S
1e�=võ�G�@��s65]B|��� \�'�~?��\	u'X�]O�Z��T���17僯�����=�A��q�A�e��[� ^Z�G���U��p���M��cx񉺘[�-���> u�3�P��Mu��k�'�"�����r��l}O�Iu\g I�2�w��%B��$��2ݥ/H@~�E�`��@3���K�͸�e_�}r#��o�����Rׯ��/��w�[��J�L~sȾ�E��x�4��z�|^�ڜ�~�1dNb��&CAtڊF#��O�d[���Wv���_~��8eL�j3�� �z�ͪ ���"�|��{gZη;�Y?)��('��VAMM�X���>���<��mkI�� )T��\S�ZBI-���6�!���vt�~W�H�V��P,H��I2jD��y��N`Q�$�f�����a�7{�:NĲC���J���x�t�
@)MT&�
G0'�C�\@�ҽ�'{��;5�~�þ���M�C�E%M(_�zR@2��>eM�9 \K��^r�o:�8	������@ﳕ&k�f�j��(� 2QY@5�Ճ��O��r������v{���]G4÷�T�A\�*d<����h��d�I�]p��oY�֛��{0�2��6���
5�v��Q�*w�S1�_���ј���<�]5��oE���r�ޔ��]?.?8BR-\��|<��<�=��������3mu�\B�ݶ�"�3���ߞ0���	�-'P}�qr�2J����|h����g%��zC�E�s=�5A����ܓR��O��I׳��r�R�������%Zϊ������/�W�8����g#Q"Q���r!�����(rqQç7�j��I�93��r-&��7�l�D�0J�JW���l���>�H�6UK�*�� ь�G��X�F��ƹ,6�4@���<���nb[ �*p+��:�����:c�._�+άu��Hq�pl��$��a�L/m����G@��o��Cm�4��"g� öF9"��ktd���M���� ��r��)�>�~|�d�����Yd{�eb�) 2�M֤�r�]sa��C��eA��D����!�`�2�R.(�����	M.������.~sF�kt��?}C�-~�2�0b��R�f���mb��`C0�N*V����ԧ����{��
!�~�Y���'�����iv�����r�9��^kW�O�y0_�Y��^�w0�U}��$ߋ�FAlQ|���_�N��͍]�P��5[������R�)hK�"�0Z�P�]��b2�?}HӶ[�M�ƐM�A+)v�� &�f˟�u�Z��d���N�����*`w���]Hs8�7R���2��.W��k�����Fr4!�s�h�1�t��L�b�S��kH\�P�0}�".*�6�K+���X@�_70��c��ç��%⼌	+Z�j��fs�D��h��Q��\d����'>�'�[�,l��ڼ�?�/���+��-�tb5�`�Q�-P�p¬�bg��X7�-�GFٔ5�B���b,��i�V���5r��}�֍iR3TXύ���%��45C����$<��O4���$��j���=9&�Z�|�?��GY*h�:����)���$zH�l�p$ᘖD;p`��[]�6QV{�:d�Ԝڤ��^LxH+/ĬM z޴)֝	!]��`:�Ál���i���Isk�o�}�[֪b�V�<rq\�>�wˣ,*�>���B�} ܇n�s�=ʼ�&��:���Ú��S�2H�ЏR�<��.eѿO������.���2>��D�lM�4%���B�s�A#��/[��1�W{̣x�L��Z�fP@��V/)i�W5���>�տeP����Dw栏u��=[YL��(V�e�r'�}������fH�uf���w��q�H%�Q�SV<8�2�7u"!G`�Z�Uk.N~Z$�6bC�O����S6�7�x��6nf?��ا�c����	�<�;�zR�q��3!��k�#$�j�Y�"x�};�Z�a�xǻxI)ʙ��JX��D��񻬣|Y�iz�X��*�K��3�[ �!A'w��@O�D�bth}��;���eqg��K�[l=�>��C锩�	�&v9��ڛ�������f5�חA#������a�u�S���MѦ�^�?_$�taN��x��I���P�t��j��P|qKjX� ��. `eK��	r��ʡnz��P˯Ԋ�h� ��-�����!w�Y�8Q���hg~)U+���v��T��KO���^܅�10�Gج���u����"1�k*r!=�y�8Ƣ�db�֗�`~�ۘ�sl��9�al��.�l���<�s���Oy/��~��呑�U�e�{:�1�����.:?��D��O&i���K�\.�ңj�D���%� ���y�uUk���i5|g��HT4�M(��p�U�x�+|j�"������ᚆ��E� s��6Ϊ��/�p�T.5+�mLhx?�\�O��'3f�f!Wת�3]������`�?K�b���ҍ+�h3�I��C���YQ ��>�z�䩜0�=C�#��%�Т^b���s�)(��l�R�E{���i�~[�3�/d��y�q4m[���ꔣM�9n=>�_2�&�hc�z��O��9���(����R(��᥯�Р�����.� ��9z:�M��[^"�����-�2�Ƈ]0j�o�~ڣ`Z��q������R���p���l��w O�j�B��� i�����OzX�-3��V`�"xJ7� 5�V/8����|��e���A��1}�Wt�sD"^gR�q�To�≲�n�k��a��Q8D�G��	�KE�酾b&֢�E.��QEiJ�D����Uе����O��J	2c�����b6]��m��c`m���D���M�/;Jd
��7#.��2��ޜPI�M�B[]@X�r�"3��d-]|H^�d�Ex^�s��\��i���tF7��M@���q�9�}�kZ��-3s� �a��vUs_��0i@��x�ͮ��w������Bʡ����թڷ�+Q����a���Q2&*sh�Q�� 3�-� Fr���p��@|B��L|\���egh�X͵h� �N��8RԊ7n<c���h�ߢѶJc�ydW��
]��F7�z��r�S��~!��̫s��X��D�>�M��-p�Ww��4�Q�$�OT�;��������RO��U2Gi,���P�=���`*hP��p�K����^�M�g`(F��CY�S�0DD$�a~=�@
K�N����$��L:��>[�[�b4d��C2��-�ƿ�����e�6ȴ\h��L���w��kr�;>u&$� .d��E���u��c?�f)ȴ�����[��A�ai��������C�7>�������uI����'l9����Y�����3�-^�!��d�f6�C����8�w��Uo��rQm���DN����lV���$���rw�Mqf4�5w@AIjo������V��Z<�?'��o��G�@)ݵ�K�\f��k���#����XV�8_;���x��77�bLO�j!=�^lf �-�hH�ꝡO���X]^�^~�
1ul��q�H���J��P���N^5��f�)b.��4��ٲ�δ�] W���5l�迓���[�����3���~C.nb����P6���3 }���kh���
�W��qб�&��W�)�I���4bL��e������C�d�AD]R�}��.pL�y�ל��5{r�u��A�G�&�*;�,�Ђ���Y���5ݘi�V�9���"�C[�>���>�L�,��S�_�����B�2M��_�:�m~�|��q~
� �����7�A�k��s���5#3��
D:�	�9Z�v�/O_y��J��G����3Gs)�t�5vO?>}��k���t��廿3,UI�y���Ĭ�)3iK8�֍�T�	͠�2����Ĩ���� �|2��~5�\ThA<�,5�f��"��El��:)*�������)'�==���l��0&�ux�},-�6|%�e`8.g�}��I�	9bnZ����N�P�i�:Nt��!��������`�����q��,�6Rǒ�\��\�  ���f�aҝU�k��"�Y�$?C��׾����x��e��^;��q�O�4���ym�I^'�WG7O�t�pO����'�2�ц��K�����������M%#������&S���@i�2�rZ������a4��މn R��d#he�t�[�K�r��zk�?�=��:�E/=K'����@Oa�}c+F\("HU�"�����c��m���QNT��#Ln؉�{gPⅻ��O�DVcϩ�'v�_+����aiNȯ��UK��u?���_i�u�u�׮ও��!��KJ4�)�#�ɍ�5x�B�������9�Ȕ�M�}Ua�4b�dīolCr	6�HN�4�G���&�y�Zz�`��0�)jA���^^6�ܶ�s�z[Nt��@�Eն�C���N������4�w�\��wŃ�/{�������}�OF�� �k�a�=�~�Tt"\�� ���=�F�L���*�k�����S�D�k�Q&�Ӱ�4o�@�5�Ԝ7��\7�*�z�g"��n" ��0�.���h�.�~9�5��R�9�o��Q�9�����9RJ�u2����5	Q��Z��¿Q�~�ǈ���j��Ȗ�"�'	x�@��d�eG�
 Ń�_�&"��)�s�c�R6\����oG���o�6I K����C�Ҝh=f�}fC��}�EUr5�����EdE��.���4ﱵP+gc������d�NF9�"Qd��c伒����{Q��4����O�
�q�i&?��Q���8$�o��M���@�ׄ��D>��;�%ES�X{�u�˳���%����U��� ��)OM�Od���n	i�P����Zc��o��T�U���r.���t������o��{�Ɏ#�X3�E]
��6��8��↔K�x5H�������t�]��4'��~���L�z�f��������f�V���b�Cjݠjzxeu�u��1"lm qL%�a��c"B��|���d�-�H���j�~I�[}�f���O��R}	MP�b�$ԣ�܍�F��a��Kp���h��^�n�.���'�$�ց�T�yan¿���]o�ņ�Y��&�0���,=0(Z���"��Wd�<�5'�4i���M����x6ބ5Y��:�і|��pL��n{i�5�:�������sq��/�^{��:�WCN`���|� ~�9�Y��K��b���%�8��n6����"�Z��Q���j�W(>���n"�d�0G�/Tږ����͑;�SPՏ����M�N���W������^K��Z�֠6�.�~���.�*q��=(\eD�h	�^=@?�tK�_)��l�J'>��,w�/��2�M?U�g3����Jǥ�5�}@��>Lə[/� �l#n�j�RK�%�Ϩ����\���u�}�w0�gY���l�i�V���K2�8��p���Y�e	V�lw��_�Go��ȳ�����1�Z���$�)J�i�D"Q�ATk�k�=���
����L�
��mE�6��:�\�"�/��=:fx�I��0���ٽ�<stvtt��ͱsw���֓�n����$~��Vx5X��^�47��*���d%���{����&j�^1i���kpԹd�Eso��S����p����8��n��L���0ov��>�>�]H}��K̩�5t6�{���-r|KR����D	������ϣ�ph���D����dh����H�Δ�(@�&�OC)�2������1�����:>h�G���V��V���q�8�7f� S����o`k������;�,F�!�3���r����Iq�
�」`nRW9f�y<����������xl/bR���"�꜐c�"*$7��s-�@�"-����2��v�L>&~!�5!��w�p�vT�u>�eb����.�荰�\�L�K�T ^M�ԧ��uQЖ�h,7����1c�ɫ��%fAs�����9������G�M(Aȷ/��l���&�Ⱥ�����i@y�<Ĉ(��'T�S��ŽK73�Rm����{�[@I�}��1#i�W �9��x����Bc�ڐM㸜��tRQ�������#rB�V�יx_�aP瀦_ڧ&�h�q�,ka��T�v=T�&�B�sy�yg-��d�E���|�����,�U��^��oFeᕂ�Ȅ�	y�s19q���g� ���
�H˩�	�u|#�s�+_"�+�0��*i7��z/b����0�-��k�N��`6zQ]J��B�T��(-c�ؾ��Ʉ
k8{6l{թ��fY�A��u/�g\d��*u�p|x?Y��ϣ�f�4�*O�&�kJ���j��O�+?+%5�f�9Lc�������Sr��Vp����'T�!{&�r����L�N�s88F���;��X�$�y��}m?�l���V Iq'(ݕ�-E�t�Q�r���AJw��B���W�^}��|$|"ɗ�B�7,�b�[#��\�1y�gLW4�����cXr�J����utaD
���n���J��*U)/�dT��U��f�|
z��j7��C�-݆ ���$���P�h��c�oYٷL�GK�x9N���J��=h����Q�|�"MJ_T)X2��U2`m.4K<!�햛hc>������2��\��@P�S���6�\(�֌�I��\��
�*��j�l����ZV��"�ܪ���|��S�3��ۮ|�")�1��֮2�Ǘ��K�a���q�٢)��%2;=X�O�U�ް[��4�E k���	'u�m��1��t��Kxm�iJ���|78h�+l��e�b������h�.W��K�Y�C�"���N�p
�I츚L����m
�&�P,�gG����y���-ΆϳA�W��C]�6�.��DW7�:��t
��.��^��	b��bB�!ʚ>� ����#�Q9�lV�D��W�د$ =�׶�!6&���FNf.�p��9����ux" 4I>�FSؗa~����~#���$[o�X**�X�B���G+�$`�����L��x�� P�
�����vؖ���$͗p��~D	k����a��I�Q�	�z`��͎�#�B�*�={���������-r砝��`�lycMCzP�40-xFA\%���Z8k.�ƕ.E;;�KmW���%*Q�V�s�pcs��u]�a�>�v
��Y?�|R@����JX�ZVڴ�W�폧`�J��L��������j���bvt"�݉�fZ6�"���%��Yz'֟>���H�"G&������s��b�zkݰą�t��k�ޝA�1�-b��Eܞ���]�TȔ�}]�f,	�D#/9���6K��b�%���Ck���IM^����*(�`l�L�k��)`��	sl�;��q�G�O�-���T��߀�s��гIhS�۝����8�SE���}�*�&�
��.i?p�.�u�l��1ַ|J;���Y��Vo�����h���U=y	�l.7�XK��
z$W�bφ�Ŕ����$׼,��XE2���o�����wE%�CP[
Ͷ]D��YO�I��qØ�\��w�5�0}�p��(�$�W���s��V�Wܑ�!�S�C0F����G��2������ C�=�[���o�N�F��q��bH����e@�@�C�����Ō��aX��x�rrrB��bF���3p����������{���vϊ\�2��n�%/�p&�m�(y�0$3i�ߵ�����q�Lј���m���K��%t{��B����kz"H=^)��s���T��J�hZ�s*�~z�^g4�Fƭ��dbRe�-7wN��E�ga��Rs��W>)�j����{Y@d��.sǷ��z�v�(�+Lϣ2����#R��`��(2���Ҵ�Y!�1�k�q�̨��_���/��q'�6��Խ+b��f2�$/���CV\x!�+c��Xs3�ޭPe�2�H���0T�W x��-*Nċ��
�J� 2�Q7��e��Q���K2\�ͯ�0��7�I�Q��wںe�R���$�H5T�C��I�~S���T���yR��S(en6��Ko�Zߙ�j Qdo�CyA�|��*�� o�9�iKWX�����u�옌9$�Uf����{�Q�l-#���n@��+�ٌ"�,�$eZt����9���n����.���u�=M;��t�ٸ=Of%�/zj e�ֲ_ڧ���x\_�s��3������)����"��GJ�S�S�/� ��Ft�|`�|хD{�?t��ZK�&���;B��V���$蹊 ����QQ0kw��t��8d>1�;տ�|q���+��m�J|��ۿ��V&�&愣�ň�T���Ų_k��Qc�?�[�C�h]�@��\�%W[GPۥ�54��ΈYD���C��_�w�FI���/ ���L�Fz��W�<�e���nFSv��{��!�K�n`�_�4e7<-�	΁�E��#�4�;[b	�`�9s�F�C�� �DE�ߝ1���7��f���w�bSӄ�48�ff0>{u7�y�ܼ�a����[�V�7:4΁������G�W�Ƣ<nq��ͼ�_±�IW(G9��L2���x�`�=9�Ϯ�K��u!�ax9��6I�S�J��Ȩ�����0:�Ż�:�O��+�ͅ�oh�W��c�Bר�nqN��� �{_ ����5-U)5�B1�
�l7��3�d���ZmV����ih��b���4�s�1�z�Qt�������Ԧ�$��gBTl.�fGB�w�	�m+'�w��~��c����q�����i���X|]�A7�^�<$	�E�d��`"v�c�CY܅t���A	qȒ�H�/|$���������3jQ$O������K yX5t�4>-���JC���8��nF�Q�B����N*�#?~�H�?�n�I;��6���"5<_Ǳ"���K�
�1 ]}: ��A���B���PWaBn%_.��Ҷ%��Ї�-9�wu0M�s>��1�GZ|Q7��`*���8iU��4���G�@��% �Sa���T���0�]�͌Yr�s�)S�Q�rk&<��3��+S5PEK�3.|�#��<ב��Uz������Z`��_`�'V���!���P�.��G�뚫��F���7�Ur�I�G�g���ykt�$��w4ϗEY(�H�
�y�coi��xD��@�/vBf(G\�V��>��HVK٬fz���1uZP�#�M0��R��F���ZL�GOH��q����)2�Lf�GG�ԩ)�v��������^=u�4�4�'�)�>�R��X�i֎ө��3�󭣻���h�� X]�A�_�Sȫ�O�=J&�/㒥���&8AJ�CM�F�l��ڶo�y5N��4}����R�����G���<��{�3��S�G3�j��WՊ�����-A��-L��j�䄕"Y�
I�	%h*
l*k4�����n����#��V�8�"��|�#�w�`�I��
cj�^T��=�A�s��p)8�bzޯW��I����Mn�CȪh�}ulV��E5t��6�;�[��d�͚Ǣ ?)�PZ�cU���|�kה�y`F䘸i�>v��%���uc]��(��
cd:z4Z����.ξ�Cvލ�D����I���U4J�v6|����T�0a��)�f���dj�0��=������7LC��I��v�6in�`Mdv��q�W0�r�s�:�4��hc�a8���Z�~e�.�!���
�8r�>� ���2�Q#%�͜1=���â8G�ĆaKO �}�ƹս���6���d�^�
m>"G(`JJ#vj�A/�M�)#9����&��Q�|Dw�cZT4qz�^&��7/߬�1����-��?+�Q��^<'~Vd;,d��Y��I�Y{�u��:�((�C�v*��֩/H�*�8=�K�o��	�4��c8�U��ﯣu7)~�aJB�R�������lf��8[;�8��fȓ�r����	��w�&	j��:;3#���sΙ�H@�a��H��hl)�m�V���;j������r�]Q��s�	�2Dz�y�ч�Ǽ���Ә0۹�$�8W��bJb��+�T�Ͱt�әU�4vdɲ1%����y�}�w�[~�QW����ȇ��p(���@��Y�KE��שtI�����YR�~��+r)#p�[g1����5Q ��L�Gu���wV=��z7*��ơ�iwJ;���G�߀D�/�_x]���)vdi	3j�}q����6t�����c�J�J�!K�����⼋3č-�:�������,�D���TAɲ<}13��I��0��"����ˤ�=ZZ��ї��sj�Qg�2}�߯���.�,l*p���埽m�H\�&͐n��D�T��%��*�0j�!�?��(�����=�����l.���V��	ȪF]���� ��"(je�=x1{�����74�A�����e�^��f}B��Tb��~�w%��4*���%�c�k��إ��x�q�	(p0� D↰����gY����6+a#K���"��l�Ԗ���I��T,�$��OT�ec�IP����[/H9�:�7$��﷘���AE%2)$��A�Ho�}y��<�r�p3�S�a^�c+D@l�lS�G�]���1����jv���N�� �,20p�ȵ�H��P2��Hx��@^o�d-��K��ή\��}W�x�u��l��������T(>;�W,ڞy��%�䵤�T��	���5K�6�(h��,Ǌe���!|s���z^3����-��Lg�2(� M�X�X5	��%�� PY"���������c���JǙҀ�n z�~
6������^]�[�`RG"�L\�W���kQo�RS*���k̆
�?����J'^HMQǅ��'%MCh�q^�n氞���8��t穃s�ЗR��u�uJ�ł��c>�ط�{{WE���]�JT��@o4���m�E�xZ�T�&�HT;�s���7������iֶ�K��������l{Q�����W:|�^�:�VI0pG,��dK>����o\r��[os�w$؍���}g "zC	8E�[	��9���w`�I���"f�7��6�l�Hc�v*6:�eH��R��+r>n���T�!�ȿ�M$/c^��<2U�V��O��u�7��'����6���V��C��WӰ�rp���wv����J��,qH�°�5�����X�� z`�7N
�ƈ>��W =�X�����+fE�"����5�T�v#����u����j�����Cd�m��0�����+�]wlv޹cE?*�ð�0<���z)���K^M��LoXLS'4��6}ζK��o�y���=�����&z��U��(]�~� Y��6:����V"0�v �	��|:A�]x��C�|�dKs-�����O&!vxc\]�񐏀*��ɳONh���J�S�F�e8�Z�t,�nR�V�)7�6 ��yyξ%��''����YZ���!~e��fPW�p硳�@�
	-�O4�XC|jF��q4m�e������j"3bqY�6�Ȏ|��{�=�LD-aL���VG�Pu�J�<O��?M��Bt1j��LiO�1A�=&�gw^�� w-�y�< F����WX��y��(/������Q;.�Q�
���X�&��7T*Ӓ��FQ�r
�:i����V�~�z��0��*~$2%��Z/�}[��ZN'��m@��&*�VUKՏ��%��])/2�Q|Y:p�{�ٻ��XW@Ŵ"+Uh���p<B\!������N��@���j�N���Җ�G��^T�8��FP�?��Ty1!g[�����AԤ¸q,Q]M���?��o�(@Z�O� �n`���r�m6�*���<B�*CN���$6����2��E	��ጳG����b�]u�p�EYvK�ȯ�P��h&!��'M��$�h~���x{]����&%B�X	T��ƞ�"*�B�	n^SB�J���+��l	���e&~�ߛ�0ͺq���9au���qM4:w�*�e�H��y�\|`ڕ�L�$����AIS��'��L V��?=K앬�gKq5q8��U`�#�WkכO�NX���ݥ��e�YAϢQ���'S+aW��?(x�%��5b�7(���U���v`߼;L1���8��5�]�"3��`��^�^�J�Z%怶�d���G|���6[���Ug���R��f����5��M1�I�*G���P�<Cߤz��Rp�qc�;88�Rs/�\�� ��*~�x�^�\�|(�":v�3�!�d��\���/�[� �Ќ=���!g�.�N����?1���Y�$O{���r�x�M����0���ӥ7��@#��Nw��P�B�8��~.~cJ�5�ߏzI� Gl*�v��qE520�<��v��9_�|(�����FM�g�1�!��@�d�R)0D�D�g%Hf�:�e���>!C;��k����������9Io�)�:�)5 ��~3�x��<[�f7�D�S���L���Nr��Kdb�	cb�y��R��px��k�_E�Q�����O��ZGg!�5�����IC��qF����,,�P�D�M4��_��B�i����A�z�.���4����Q�f*b<�/�Ws��!�Z0p�����Z����냰��^͇�GP4*�����}2�l�;�Z�Ԃ��WL�]#��'����"��g�h�y�y��� �(� �E��%F'�my-z�R2�ʻ�WsM�x���t��_��OP���;6���F�������ĉ�kD	 �t�ZR�)�5�Q�������pd+p�wy��j.*8jC�ԥ��̮��f-A���Ji�Ÿ�m�c.=�x�!l�-���W�����/����跾t}��\�g>���r�ژ�
��K�u���m�U��9�|�.��X�G4�ڑo�G'�s�rt��X�s[��� ���z���Y�����jɥ�p���@�?jd7��j,�9xڮw�%�VQ��6�Ú�L�	�x�Y3�o~�U�̪C����ꪀT��4��˺�dlZ>7&o�a��ǔ�T2�$a3��[Uw` �۠�~Z���0R�+�{G\��c��Yg��٘j�<AE��pwa���J��uY\� {��%S���#U-��d��W.�\v�F>�N��ܸ[edӸ��{�`?&������_�Bgq�t��Q�E�e�"m��i.9u w�gw��\%Ѱ$O\�[\z��$#/�"�*uk�ď��nH�����&��]�Z���q�Vf�:�l���"
��=i�R���w�2���>Y.��M�P�v�b��ͅ��z'A�����OY�l�6�΢kY�7H���Wꝇ��F��Qd�T�ɞZ�T���^i��ʼC��WL�'Q�[��K��v�;޵i2P�GX�����eKKt殇:���gu\�Ѧ�?7�w@�iscLζ����O�����<�Y2�fQ��;��e%��n[�_sڬ�]x1�	����- �A�5"��FB��*~���0�3�Br���G@� S���,M%��׸�H�r��~�ԇ�޾�+j2ߙ'qp?�F��\���H<5�h����5��QǨ*�Y��٫�u��ىlP�TlM.��Ҟ�.��w��<2�v;~�L����r�=��'ռOz5��qO��	x�e7%8���`u��E)� |�驷J	��B��ˌc�q4�a�1t�W�&*�����K9����`��P�����N�����܄����hT���G�@O��s�/����7����!��,���i�+GM�Q��A��<�;ey�C��]��8Bm�i��\��
�qa3[5)�Ś��w2�(�~�ٸ�zdǆ�I��s��z�<Ϸ =��-.=�eM�/HR��7�@�C�$7��y�2�h�B�m� I��*Ie�����������5a	[�<z7����ڞb��	dX<�	��=ۿT���Ji�*KGz�Ե#�t'�e1bA��}?L�����{���ț�#�J���F���H(�z�<Ͽo�`�'��6~e.P��R�;Eq+�|������M�YQS�;��z��zf�tz�j�� )�AO�|J�5�_j��xEzU�kFG�]���F�~��,4������Љ�T,X2z�/��{����'{H叵���g`�q�EG)�y�Y����C��Ҽ������e��{'hj���\b����>������~����t,ȏ��	p�~����׾Ko��a��Ρ�!�T@��t��k�_�����9�=�Y��J3<�R���E@���'�)<+�oBQ��l�[����g��}[Gv�'���
<���5Ò�Ԛ�>����M��R��mgW~ ���i�]����8С���l�B	=���0ȉ"Q����I=�"��1����`�W�5b��M/����! g�U�� [��e/�	b`u�g�Ӕ��`K<*�叞��;��@�"b�D���j��l2���uM�L��l��s�{|�����G�,�5��,��n�q�Aj��%�6�Q�;rr}CӮ��	j�Y��^��i�kH�92*w�|+>�X����j<|�����<���xA4��3�n���+g��׃���J��4b0�F
jot�;^�^�o^��+*
��dMpe��h�aUK�H�S��'"�6S��WB0o	���-�fD��%ry�']*�Na2���!��^���!�fj�ò�� .�8tz������FO��;�������<�R2=��D���/�l��u�����&�Ѷ>z�&M�	w��fM���r?>!���#�G����v;0�UE��#��Smˆ�$�����LUY�ON�Y��ץ��ij��)�m����^ؽ�5_�6E=���'��~��Ĉh�q�x�p2�,�hY3�WS�d ш��J�(�Uq�94���  F�WZF\r��\���I��3�B�� "$B��'���+����Z��Z�vh��<Pf�'�(a����Wj������(�����9�<f������c�t��8L�5%�gc���f |�E�>�z�`9xď��vB�b�O�̼"�䦞����C�DI�_�~[��5��7��/@S�c	[����{D� Cъ���bEZ�]K��������� zDA��:�N&m�ԗ�]D���׬;���Ge_�=T�U�=�?}{��6�A��E��pL�Ly��>E���ϴ)�D��H8�L�E̶��V/�'��7�����{��`W�$�eC����Ҫ�Rp^cn��mJ����o�V�&�8�c�Y1p���z����*ۼRnÛhl>��%E+�#E��o�#�2p�}�4�/��69�6�h��mᏔN{�/qh�<6�M��p�hk����XC/�f�[�@�P4'�Nfk5�b�sf"T�&�c�c΢�U);��W���Y�*x��N��1�W�2?�H�-���?�[2=*S�1'"���s�Y-S;f؃r��N���r�;�I0�vL��\rd�����V�Klӫf�hy�u��YT����N!�'�R#V1�=�Qצ�@�8_�B�D��'W\m����%>�y����-O2�zZ�FT!bv٫g4�陹E�ݎ<�o.���@����O����mo��O� �ng�����$��xu;�H�XxA�S������|����c�|���#�!�T?�o�R�s���B��2>�ԇFԭ6��:��~���e9M�yf��բ��8�R�L!�����X�Ta>܊S�F5�a_�Qѷ����F|���!��.��w�]�%�>|BƁ5�Lt���×��߰CB��w�S�"/�f���<��0�gп���ܘ �z��QrWe�-��Hܗw�>/x�Ϭ�<S�z���n���]$Å���N[�k�XoC�y4��h�d�|b7�Tq �\��.1Fw9���Z�HŻ#CQ�{�.K��{��6R�-�7C�j�c�X�=���&�oM/���^.�-\d0���1 ��IbO�m3���[��~�Ve:a��(+-ᤪ���i���;���v��=t������v!�~�8��k!��,�{6q�q�s �I����M�?���V\RI
��'f�=`�"�1
,Oa��"��T9��-m�4N�TJzT�n`�E�Y�χ+ҕԡO_�ُ�|��:��$0f	��X`2��)�ЅA�F
��q�kɴHy8o���_2��G�,[Ӥ�<f��A�^k������s7�9NN��j��s��֌j��3��l�7Y4��+O3qD&���y�&^�N�A%�/�J�&��5IC�\<ӌ�?cU�g
��{1/���py���P��x�,��}�j�ƬXIZ��d7_�I?���'���h��Y��&�L �d3��LF/@׊qO
kZ;'iUT�_Bb��I���MR�\��&��H]@\M]f%���S���.�DyF+B���)!�	�OLb��{R��d�5,�=�P�
`;�����
�wZX���W�i���[[e<�~a��"\��q�=�O�ӝ5l�+1��'O1L�`F����6i�����<.��6$��R�ԗ
"��^��HΝ;ؼ���v�DT�)~	�y2wO	4?�X�#�yR���Sq�ҍ������E�֑l�K��`f�j��2�L�W|�%Vk?�l�6��A�U��X��6V��������F���~K���w��s������Q�����!�C3g)�.��� ��U����#eO��i�0!M����L�#�ˌ�S 47tk�^� "�ⱇ\�M�&O���1Z�\4J9��12���F�-`8��3��Y���8����0� �µڶv���#RE�x H��?�c�V����
���j�k�y�z��~��y��������Ն��B|��ư��_��%;K��A�l��+ܤu�2�1�x6a�48n{��	�Y��cK\��*Tm�$U�;j=σk�x��P�OOH�%�m���%�P�0/&�9s�q�^�B`�K�<y�('nf.�FR0В����TÒr����=f����g*��эΜ1V�C�}3	8WUA�T�q��H�YWF�����A�>A���m
�t�1'Ϝ'�����71HD�
y�@�p��m��/>q#d��!#����ƥ�\>�1e�b$��{��$����w\@9'o7Y_�K'�����vh-�}�w��6��ԃ���@���_�R9��?��;EЙ	q����N|�V�&T��`�0��(���� |~�#���������"�3���+���H`��$uE��=�Tj��q�A�t9|{��y�Q�s� ��R��غg�}^�K�=�
�n ��,�HS�5j���B��M���	���'@�4x`����E�ڥ��Q^I�ܙ�_�=>�7��-iծ#����ׯ!-�$�W!���+R�$݊$�a���EvA�7�4R��f�V�d�����D���`�S��s؄RNժ�ⳅr����̤����>����1h1ju����MJ�@%_7�3�g��i*����7��`���Iy�9=c��V��k��J���m���^wkm�ǡ(�Q���/�,p kO����#�0���h��%u����x#��@Sl��met{C���9�^=)Ƈ��}yj��SnmT0݇e2,|�%�~�?�/��q��ΞI�0v@��`;$�){Ni��ܗ��E��P]-���|�X�ta<3�Ӄ�[�V�I�#%����ٳ����ieO1���T���1����8���z�S�f�!������͡���[
1q1^1����1�T?�%貗�n����%S�oM<�RG���5� 咯ʘ���s���g�϶�:mֿ��Z�quPb��Ut}"DD|��p;��ջ��c��)�5�kڱV||7��&�/D��ޔG\��M�������f�SM��޲�0�[>D�D_��Q1F��4^B�y���*	t=�V�� ���p̳{���>�zV�_̟��S��6�^��H���ݐ�~Z��e�g��m��",����7�Z�;7�'9��~�rͻ�ڂe ���V���+r S�KU��v�?�$��ʶx�&7������n�X�}Zॣ�#%2IW��Pެl|sm;-�a.�P�[�C�\v�k0��bZ�f�h���Ҧ#�� _$��8u�C�G���0ӯE
�!�?�#�K��j�E�xXNa�ɋ;�V�T�w��S_���M�+m0k3�����K[ =�$狰��S^�9�]�>	�z}YjA�������L+ f�A �O@e�7f�^�1��b~�*{<y
q�_x�j
]jS����-j��W��6����*�v;,��� =�lb�bA3x>	2U6A!f��U��HT�pO��Dw`^�W����o
��6��\�O_���Y��ן��	�╗���ݒ��Ò�:z4�_�Z�.�F���He�2</�y�D�kfb�>r���@%A[�L`+��}�J�X̉�'(�ID�5S,t/�g�5 #r[�зȑn�a䵝�箁� �8b��#Dt:�Bx��4�����X��;�q��^�		��+C�o��Hs��91L,h���GZy���S�A�Q+�6�)Nd^ZW�L,+��,3���Rj�Y�p�M[��M"ChB�S��k՘_���t�j4��_���b77T|�B���}�<�E�6+��h�O�������gl�E�e&c�n��0�����p��?"PL���*ow��&��1x�%���ï4�������I7g���nS\ޜ'���(������	��@��� � ��+��Mx�W��?&��i����woަi���.���� !�����H���!KH8��D�S�G>S�g�ܒ�>�k޵l�X���rc�{��n���	�´R������I`��4�!6�w���Ol��r��k�+�nh.:�d����5E.�C4a7u���.�'����&��T�N���h?��hS���^܌_�Bg6�TkLl�΋�܎2OZ�>�X��Mxc5�o��R�PM�|�HQ]2�|��ƠY�߼�0%��b<%I��D��=��E8b�9�.���^���ׄ�H��:��%��t��rZ����R�BD}雽))M
}<�Y��ۇ^�wP n�!��'��m��7D�z���V������M��'�����!t~�x��x��E|���w�j����L�3ߙ�y|�'��n"�*t� ���]��ʤA�)�����B�	?�vՔ�G�y6���p�:�����̪�-�JzGT�q�����C��I{9�+�<Z������Ec��A� �:7{��$��&�ހ��u}�U�Q~�Ҝ�Z�}}�M͠pe6_h�6��13�h���&�ӋDW��j�-�����G6�9�