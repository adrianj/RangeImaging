��/  �Xt�`$�����My<~}�A��5@%z7�FH\�0��-�9EMx*1�s���v�G���n�2uO#)�Y>�P[!W�n)6����o�hY[�ܾʰ��)�q�3����ϺeK�^)p��Hz�{%,rU���_��^�^ۜ���l��1An"3�"�����o��LV�laD=tp8FΡ��'�N$4b<9^���_.x.�S�}��_�wd�rV9Mz	kb�X]!��:J�#�7�{r��x���:ό���Ȱ�2y/r��m�\�R$�<�V�1Y ��\?;W^|�bAj������h�W<j4�U�e�c�ދ�c�k�1�xix�`J�_f�2�	�ӊ�Y�������-�#����R�9]#�G�QӠ��
�N�< ��/F�+*��?<��i�/����b���X*�ꂖ���c �c����Ҭ�rsoEAC�XZ�M[��������}21�N/'S�2��b� eM�x��44�hVk�
����*6	���ҡ���㛜�
��>�VCޗ��9@�ܴM~�����~���:�[>�!����W	)T�F³�.�sA�Z��R�a����F��S:YB0:�;��Ť��27Xaϙ*);���%r�(!d5cbj�!/Tל'�N�!�w5��f�_ࢇHڊ�U���W�q��)����b"���bM��T��m����7~�.�<!�o�0��`�ˎT�˼�c���&��;��Ў��<���ƞ��s��X�r�Y�����/a>��_�w����9i�#\����h�c0�b�\]Θ�%`�@] �:s���m�d��Z�s����F�f͜��p&GqC����ι�L|�P^L�&!Aw��x�9U\�+�f;�jI�(��� 4W9Lru?�F��'a������N~���B@M��bf�9I"ei�j�ySe��r�o��g��qP��&p��M�����(qK����4;B�y�>׮��f}T�"�|��f�
G��՗$��`p��Z.��T�F\4��hD���x��O������ū��D�'�N(cQR@M����饷���a&��3����~�~V]�"N����{O.���ת<}�pgU��Y[bЍϠ�g�_�̿��&�WA��܄�Rv���c� ���0t֛ӄ@��2ʅ1�AR�t�@�g�,dP�w-�"����5� ŷ�u ��ш�AF�|�:(�T�{�P/	��a����VJ몢n❬�_d�3� F��x��0�b3� r�q�]"If�Q�L��N��za��������x�E��yn���;�֙��P�� q�a��h�"oI�����>"4�e�4�)�+�{�ǉ3�\�<T_�D�&�5�����^����9i��{�"�f(Ub��`�{��`&��q�/���1%�IHzAUz����n��C�/8;��@8��x>�C��W��g��a2��%H�b븀�8lw����3k��EH�Vg��~�1��ٕҐԻCk9���_k�.J��I˼PCO��Ǥ�5���e�9ψ�Idw�)	xDA��T��*��\X_�^�2������0`,�?"?��'4s��^�{�H����(*{5��UBf�x�8��L�]V ��GbzE�!��A��YR_��ʓ&����jJ�E=��O��S^j.Xw��xz�`M����:v�B:@W륪(��O?�������N�85��~�G,�hGC�s���"}Y�J�p����h M���/�3-������c.��� /�{#�"�U�VҖm8�8� 9�_;뢿�A)��7���u$�p��UP�VR�IK�S����܇47���2~����)��XtU�+��6ud��`��s�n+�եp����
����Z�F�j�(sW�tv��g:�ZgIפ�+���u�կ)������8��2���xo��h
6�K�F����1%�[� ����u�*h����x6_\u&A!���U�c`��j�a��)M�DBϯ��A�9X{2SQ,����	왑�Hj#���Oǉ�c=m�>��l�����H��V�D�x�ȿ��(E�!v×(u��Yx<|�h��g.ʪcr66�S�[��:����������W��hﶍ.|�2�6	SY�.U�y,��R`ֹoM�dg��=[�WJʫ��1��u���FqGr='�>�����[�a��[퐹6⼹Y��N�sc��$���*8�`�9��@���8E�bh��EA.�{$��9�bˮ�u��XJ|E�f��I�`^�#NƬ��� K�aہ�@�g�{�;Oێ,��zql��$���e5,021�OU:'VH�:)=��^�v.\�UhL�]���2���7��[�D�;֥#���we��s ��Uv��n���є�|�TC�
]N�$�����~B�b�*�{���v��E��߲�z��t��8'4�D랬:�<�H�^��k�~Ml6�Ɉ �������=���x`��Y�����Y��{$�i��V1X�Jx18���Y�6
�sv�5�B�n�p���<�⼽;�%�;�>\��B|�3��)�}�$�V����i�q��p�>#)`�v���%�/YE�*�8�P�!ڷ����H�:YlK�c�j�P��
!y���^�j�ơE�D��+3��#I=�U	g�� �=�#c�L5+��8i��@ Q�t�P��DE�`�j�ɷU�]QQ����Hl���x�j�ӃWɀZn1=(��t��agq(��?�!���/;mj?�V�8�	'>�XJꞹī� ���>�ddh����U���)q�`f]mD,�y�T �D����u�u���]��9���e��?�^E����7R�3���8������l~�G{��f���_��/����*i*���o<���� �C@�ЖM%
}� �N ����;}�@����s�n+b�A�ׄ_*(.�`JOق���Ph��d��%9n.����u5�5S�3x�D�����9�V1�"X�[|�C�s�H�����[�+;`o����K�V�b�K�]_��1)f�;>!���LeH�,R��6����#V�<��;�Z���<����q���;8#��[kU���U$ܐ��) ��I��^(�X�ZjIݩ:�M��՟p��Sr/��+�I����JC��?�9�Z2p�8��E�E���Pl�9/�{��\hDG���=-(#}���`�"E��UB���pO?�Z%�U�DW#X:����ڂ�D�����j�64��l���Ŵ�k�Yt��a>��^!뇲�7ɩ���C��@KC2����7���|Ow�Xc��ۘwaW((k�\��+_3�W��a�]!G�Qm�OSׁ�i�����t���/\�M�R��m�Є-�gf8�u�"ǆań3�٬LG+r��GK�g��*��x��"�I��<g���V�H�Rc�q���	ԖR�y�����Y��]�q��//����x����<ľM{�m�\�o�s�_�Y�4��r �I���T<d�9D=`����E��v/�T�%��z��<Yе�S���R��j �h�_����^��:+��2��+�u8��XsgG����y���yՉ�{t��o1ԗcg@��4�����a��h��&�k�\ �@p�ZH�͹�4��0�$�U� �(}m{ʶ�"k��Wj�T�J&%r���w����\� 
|\�y�
����g'p��n5��1Y����#_%�t\_gi%��"1(	x5b����4�M�ZVxo_Z����_�c�>&�%�͗-�_����:�d'��8���8�@\yʃb��ѐ����+�۫�O�븧�f����k��BED�m�&���$�s��AȰ�&ۜ.ϰ.?mǡ�'��6|�?�8���]�KI|�^`��V�f��@>i�.��7ߛɰ	��S�qbz��Re�<w]����8Ӈ2Ŭd���e�'��?u�ko��Z�)
|����
���p������5�'��8�j���R����'���i���9�k�}���O���WfV� P��J8R��Ji|�/�@�ܰN��Ͱ�֏F�F�����Hh�1p���<��]�������.r�i���O���#�6/W��8��%k�d�F��ao���R���w�!u�Q3Qh���ß���f�4k��i���� �&��F�����X����%Ś��%:(�*1�e�D�V����bA�̴�;�T���v� ��z�^e|�I&"��|QU�zl����j�`�W��7����ґf�Br^k�w�%�)8�x���� �R{���� 0?�S.<�eQL�i'e���>D�s-����bnj%��ê��̬����j���ө���G��ouk����.@��1�����QK���n��{�<v5L�e$(K�L/����b��X$��%t{+h��y��V�/�m
.ɤ�S����[nA��Ib�x��ʫ�%d-��C��:��8�8����Ȃ�]��G7�o�)I�CMy��B�\��rp�ӢEped��U����o�)H��P��!�!�Ui�ݘS��5��#/�Ϗ4���t{�^4y~��MO�|�^~�G�R�t��>�/��!��it=�ۙ���t�M����b�^楡*{���r���g����b7l}��*�s�7��6~�;��̍6�+0.����X)0h�2j��]��eo�U�I_�|��Je��1� N�U����:.�t�s�]#m:t���~0��^����]ѥ�j�QE[�z;�,T��HX��I����8���3���sX)q����:��Ւ�O�����x�K�W桦���4�k��K��m�2����;�1�=�H]�c����(. a��^��z�zob؊�0;�&���?!�zvL�Na�7���/[�>y��Kyi��ޡ�z2�*�b�{4����7mNc�!�[�$#mk+^u�|���y��Q��m|
���˫�HI�<y�{-M���vp���B���a�8��'0u����<77���/N4����$}�#�}~ȕ؃ȔC"�F�����o���
#8��C��k� �tc#��&!Ks:�I�Nh��Y�/�P���N�AҗL�⺳}�e�t��,+4��8��n| XRW�M<�I\I�s4pC��3#�C1��?��޽)��-�J�!w�����d1烈� �����@�׼����Ȝ�8[��? �B���K���peɲ^@�j=eb�5�t� �|��t�`,�*�9
��Q��B�|��}�J
%� |PnV�*&X���Ϸ���jB�&9����F)�c��޵�O�bk�A��\��S��rR����=[\����J������x^�$�>��)�?��Ƞ��6'}��Ԑib*K*�M���fv3|���|ʭ��͝B<�j�#�@ ,�7<��4�z5�uѭM��@�ת?�p�J�B����!��z�1�1�;CF�gD�3X�6s��p;�˭��cG{aY��]1�==�jT���JJI#��ϩ��1w	oGh���ᖜd/����M�4��p~K�MGъB��h���
I h̍�|�vB����oA���6�}?������!��,��嘫�E`�M7��ʱ��.�ހ@��V�u��)���u�c��6h��]��#���u�k���0x(�\A2�XU@*�������GK��EN��_�Դ�W���������w��Z�j��r!���x8�$��}���L�KA��R�KUk4?�puED#��i�3k�1j�ॐ��������i�-����H�����{�j�Q]��覨'}.%P�T^�͝����(s�.M���x����4֊��k0`����Id��ɘ���Q˒���O�^�ȧN���xI-�H(gPµ�R2�f�N��<���Zh�|� �ӹ��DL��3*�
��)��$�h���1?�P�(�W���::��\�%����:1݌3�C���`?�-�����I�>^��/��6<t�r�T.i>�:k�tȵs��Jk�@+�ˑ����R��L��"��V��Q��"�1�d��Q���"Y�	Zv��T.�{([�z��4`��Ku:]�5����/ �������t���(�i^�N��f#��.kg������������qpF�3���'�.�or�b���T	��;��������qU�?bG�}�𜰺mo*u26�Q�eu�rC�L&����GTٟv_ɝ�5)��RԷ�P?K.� T���S���z��7��ko��\ś�7�sW��}�J��;�bb�1\?���@R�
kj{�i�hKĈ����i�6��z�٪�5 kH���.e����cی,�lS_Y8��Pʟ{�.�bc�-c-���Ep�
!�-�|R^�����b\sMm��?�v�h9�
��t��u����2}�=���y�]�	��@˦�Ĳb
m�2���XR6��q���mĄ:�.���|�B�W<�c>����6�c;�o��ƵTo=�2��:6V�T�H�*�(����'p��FѴ��!]x�L�
�O"���y7�r�5x���AD��%N��\f���'Ns��c/\�.��tΰo����H9�U�f	��`',�I�:�J҉"B~�������P5������R��v̞d.i-��sM�0Za\����K��W��q?S��:��Ʃ�}^��Te�~��Z��w��3���Vy����K�?%�`A���#c�6�0��w���hQ-bU��q6��n��U�~�����z���CjO@t�2S���[�ޫ��ZLF��V�'�B`�$˻���$��o3;�T�!�"l�M�U��`�{n�y�E��A�sA7n��Ԇ�8�'��g��0hŞ�i�aU׼WWN�>j���>���uRyi��5�q�8�J�
�b9��[��z�
{�6bϿZ�i�zl��h�9Yoث��Ębɑ�_��+�<�=ȁt� �<lL������S0�ŵ��j� m8e/�ul�����QC��Pj6�{� ���z�'���H�H&Mv���۪�C��"�T�ėݽb�bB�	|N8��;w-��?�)�;�7����`��lu"��P�z��C	e�i{����߬}����)�ͲD���oÓs��K\��e��3��<~��K����%4��LeJ�T��_J�FzO�Q���{3�4�$*�8]z�����n�gid��d�<��*N�ef��_�!4�,��vCy�s~W��%MR4�7_^&a���s��ƽ'#�\
)��/��m3��ǒq"��=�`uBq�4g[�L�-O�����Oc�7ߧ�	��+��t�j���=�
]a��]�Ζ3�r���X#���Ѭ��]�˫Rz:��}X;{'�U�Z��R�Jy���q�F=��$�9��./��Y�'�RY�o%\�����5�����4y���)���@���gI/�Xc�J��$iG_�kb)4}|0�)��S�`�$!�[vv%�E���ҝ� x�]{�����*&=ˇ�:��`��T\S�S�{���o#Kʉ�]�v��a�B �ך�/��` ��ɕx��D�g1я����8\P�V�������6Bx2����D�0/��u /���������.G����N�
�%�n��Š#\�}�
T�);L���s6f���&]����V[����r��C�z�{��_��jA�83`��z>wE3pdh�Z~�C �.�q���ʡ�#�j�� ����}����m#U�e��.�f�op�<���͗���_���܌&�&?�����-�&�bb�gs,�@7{@�:��q�I�
��~&Z8��{�Op��/ɡ�h��4��Lu
��m�l�;������"�SV�K��J�x���N��&���虇}����$��!��C���?�Cmi��P6U��� �~* 0$bE��1�Jt�Aw��R�2�^-{g>�&<s3���Iq��X4��jS�He����������{���@x��z�Tu�����ۀ}��7��
Eìe(��<�����^����[}�Y;Ӊ��)$�^���z�\�����`S�щ }���-}�����᜚�lk-�cYpk�W���l�Ռ�U��
�n�YV��ւg�-�V����K�����%8[����>�4�v��`B<A�\B�[Q����b�������Ù��z��"8�v/��e2�p�C֜����ų�FV�^G$��F
O<�,�NFj��g&?�Ԭ��n�l�$o�X��w�^A&]���y
�Ⱦ�J,��*K�~�Bѹ�G�d���%� ���a~F����]t��2�	2����|����@����#��v2o��k���2��W�� x�+�����w�}?M�=�-��X��Y���ç� Ӄ7L�+?R����w��N�*�ϪC��R͙�l�r+6� �f�}~�UƣuK�E�fO�}���KV����(�7���j1�W���݂��e�����r����ۊ������.��k�Ӊ�L#�wE.�%)��@c��b�H�2�AM�[���g�E{3���ɹ�!��t��v9���O���P3=?�7��5ʅ[b��l�0<C���5�g��ҞJ:������/��� !�������*� yk69��֛Qd9�cy�*6ٜ�O�Xdx��)��ᬃB3�=j�q�5	>��$��ڒ���\+��9:(}�?'˦R�^r��Y@3�����}n<m�
w��	� Ӱ��T����J�R)	���5\ޯEf�ee�3|����J�0�u���H�|f�H5\|���v�N&�r�4ṵ;�Hȕ* dF���iN�_��i�ڳ����tv�L9�+ќ��lp��ًZ�G{&[3*��=��&�� ��OI�Y%�xN�k|�.��_��KC1��X��_�A��q���dP��j��K�!H'J*�lh dc�1YE��+`��laL�{|vx��[�Z���3�i@�"V�\~���G��ˤ-:���P��'MP�`3,GY���n�9���Cl�Wl��%�p�yw��9�.�o8T�$��1Ԯ��\}�T���uF����&906T+.�B�3O�؄yzC�-bn��=�dQ2���RUZj���c�q��&�^���
Ѩx1>�r��߈�޵-����"�m�Y�N�t��N�1��:}��k,�/=�Yi�I���bȵ�E/��yB�Y����?�c�Kd��,�9�{oIS���!�y���4/u�PZt�q��~?�kB�'b|����Ǫ`YZ���+K	�
���6L�R�_yh�i�����!^��b>�����]\���(_i��|��CZ-�/�N̕��S�n��0tR[��F!��2�H}��r^��I�Od��?r3bOԶ�.��<��;�k�m8&�
�M��~�������@�/���.��3fa��2�eD�����/ד���oW�"	���+�,� �5�z�����|<�*8��?��a5�>T6i���C�K_�os�k�TZϬ. �{��y���+6��,̑���j��l�5��ĨWM��}��^=щ`�,�Jf�2inkw˳��Ƒ��;K�������%����	�Z��4U.S����+?&�t��t�c��~�k�0``h._��1.}�Y�j��4~�{�?���Y|R�r�Z;Ao����Z�� �ߍ�d���d����pi154?̥��w����bkwٻ�w��Ⱦ�X�����|�S����Ѐ���I�P>�*�e��y���0MOy��30zz�]J�'T��w��
��> ��$�������KLV���^���f�i����jf��9S�O�I�-��������ծ�jn�Lxc9������e�����K���Jʬ��
IT�_�}T�kC[�E�j6�4#��B>S��-�5��=V-v�}�{�A%=:�j$ٵ�t�q�����^�T�X�o�rw���(@!]�1v�3_��QI�3�+��5��G|lL��-xö
��j�n�2�+_A�%=zz��٩��l�����o�\�7�Y�4��=�NC�(_s�7��I���K���V�3���w�g�ԡo!�*��)�X���E�-�l�7w�P*���)���S$��,�NJ7���������`|FCcGJ�i�GZK������~����b���̫:b]�D$dn��2.'�pG�{��CRp�#>�'���iՆ�;a}u~g�Fԩ�{�H	y��鿎L�_�]����^P��˴K��\3��V�7氊�I�;ǧ�4��+���j��	��%�	�w	���8���g�Cm�X�r����	r"Ax�S�)Z�Hp���9	�r��T�93<aw*��������$�D���^�~l��Ѯ*\�hQ�y���J��9���,\տ]���Mzf��J�Q�5q��Ӎ�A��nm����֓#�?*N�9�F�6!��mW�ZͰ#��*YnjQj�m݀^m��=p�r�h���m`�5�g����Hk#��݅���i��r �ء@Kên��֣�>In2R���!�%��ῤ�=�¼V�%M�a��������ބ��u�L�N��(s�9Q��.��O�iL*������.��#{���t���ā�����R�Y	G@���.Q����8�u�[A��,84��G:�*(++��,�¸�E�L�X,�t^�oe����$��ˈ0�-�I�~�w�5�oШ�ޣ&�y��$�sa�W�tL�OyPT�mU����]^�tN	�b�;)�4�u��k�~�D|Hl�������,����dK��{�&>�z��(2������&�e
"p8$�6xh2)�ٴ/ON/P@ok�ǃ���Pǐ��Ta�S?WX���%@��`s}I�4���)�לKZq�.��j�h].?���	�e��"��_����U^n/���\�2���D�^�w��!g ���pN� �\�Ĵ׵�fwMvɂ�s+�/1�C$2�4��J�x���E�?4�\~�*�,;�2��R��B��)-@>t���,}�}�5��Kע�L���i�a�bq:Ƕ�%���!9��ܲ{R>?ss���j�&�9�r7i������/Yz��5k|rMXU�O�9;W�����`��&�8����wǟ%�^�d5���_�ͯ�oUv��"s�� �,S� Z�D8q�V@B<_���Q��鱽Pv�ɠ�jbAL�Xg�`r�+
3#��/1�{]��HS�%9�.et"�����𧓫?�i1.[�2���?����?MqZ��j�`�;���*'�K����$)D ���|���Q���$�4_��ͅ�#�M���V�z���c)���Q���ųo���1�	[�E�X��"ͤ����"���C`"�H�w�RS��5A/"�<�퇖������g��Po�ႭY�0�C��'�.Ѐf�ks�޸�փ
p���3�Oj�_�yXB �EX|���O�j��h�6�0�vϹ���;��'kY���������,��#P��7����}��� ߿�ŎtWT."���K�gW�,�ez�>��ϯ���� ���� ٩�C�3�yko��z�c�&(�쉻��'w�4N�wo ,��ƭ�h�C��旛C%����/|MN�q�=�N��� �=���NK��VE�1�9cڽu��و��վi�z�R�6���+��g5f�ۃ8�����J��Ï$$~����`I���ϱ���T����>�/k�3����:2�v��FS�����\����z�ސ�>&.���/q��h�n���}�O��R*��2C���t��@�cتuH�VOebǙ+�;�3u�y?OaY3Et|��u���nʉ�/�QBIٖ�]8Z�۴ �UuO�2�7��Q�d��:�w�������$���]��<o?Qw���@���)op� B���4��KN�ڦ�@���+��E�1�f���A�F^A��x���󕞄����+�A�v۲���|��Gtu�n.����S�&۸*SdG>��47�j���������_v�N�3��-�:gp����v^�t���&��XaO���"6J%�-p8ڀN��Jհ�]��rb��B�j���Y�B2�!Q�N�=Y���tΜ����i-Ic�m�?ۆs�qO9�Aϩ��/�K:{�@%)@��1�zp�@������ȷ==@��TMuS�b��8!��0%Q�Z^��EC�SH�xAeM��A@-M�}�W�o�X��sǇX,��$��j��Lo/�s�̝�u�=a!扖K0i��;�Z����,jZ6����_����M)�xO�!#>�؊!�r�u���=�D��v@�*<0\c[@X�j6̪J�.�yĸ��]j�p�KDq�#%M�8߯�I��/�>%H?O{R�f�S��/+xF��\uR��E*��&МQޔxk�,�-�շC<���L;���F�g���I�����R8�!l����:�S�W�Ƣ����`f�R<N{b�E~_E���� ��. �?��3xW=��ڈ"$�����
˶괟M��Ѕ�����P}[@�PP2��3��(��]���ș"n�sC�h���>W�J�J<�J�Ʋfс��ڦ�O�)j�/��Z����w V�H�x_����$�hR�UBM��$�.ݦ�W���^�̧��G^�����3�cyq�
�5�YQ�C3]~��=��̝�����L�������8�H����Z�����Xf��o��L���O���w��<l�6f�4��r�!���ط�/�׆��TE埔����h�YbGĮ��6�^<5A��������m��?��w�J0Oa�������%G*T$�\fa�'m�T����}�tn��&�_8�z� �������L�P0��������f�ϡ���I��X%��{R-�L���t5k��_L!j�3�ԇf��Ѷ�L��.yd�yM�ƁѾL�
���J��:��*��\ DRO��u�k䊔D^gAiU�쭳����4��jZ�B���J�f�&��ޜ��[��ⴒ~�»����%�?I�χ벚�'*"����Ka��Tn��L���%�D����3 �dc-F~m4�j�,�	m'xXc��#	��j�EV��*��H�|�����(&�x��u�3ٻ����`涯,�9		����N8�)����=���OK,�!c}�� 	h��)��t ����r���r��Ь����UrP3��)���M��*�5�3?5�h�K�LЉ�SE_���k��V��b4�~�l���c0�h�BaXӗ�Ȓ$��tS�qA4�R;+�zoՠV�h��&{ ���U�q�2�8ȸu��'r2���5��wXVn;=������+s����+/�-_��V=(��ж��gJ=%$�;�*����V�N�[�C�	�ܜHs��w4�~���:�u��E���1�5�C�9	��N��Aq��l��k��ߩ_�r����1��nS6:�~� j��5�{wH�.�����5�2�jM�;ݴٜ	z�,o���/��D������4,��X̀��x�ف��Q?o*��1���z�r/�^2��z��AEFA�����O�,�:4d�D	Js��0�V�}W�jX�LJ��퀔V|��LO'a��W�'���V��͖xUL�Oa�*�4�eժn��`)�z�L�F����]A�H�y�9���:Jg�:'�����C�JWl8@��X��l@�f>q@��|j;'s��b�	��J'�	�*W�F�r�~ԢfܸP;^FI�Gn�à��S��/9��G��8������l1j�wv�Cv#�@�+�{�2��T�ٞ��9�,�Z����P#�����V�����[
Lg`��z�C������G@ o�%u�T��\�>2f�����Hz�U��P1T���Q��;��RA�@l���Rm��j&����*iAm�W�C0ۦG�x�Q� ��-��o-Ǎ�ԏ������n�ª�7�r�>��ս�c�l`Y�����@�7b�9%�F��;��C0��iIp��G��N*׹L��G�7�l��`K㊲���e���Xa��J�f�	��\B�뼞�k2��}�f����Vy�]�F5��:�ϳ�p~]����0J���LZ�S��]���P?d�d�+��~!ftI�v����E9H-R����bR�49�x�X�0�uzJm1vZJ��b)�&vet�u�/KHn{�̜ؼ��l�j,M5�1+"Rz�ά�"�@�����4���C�X�����QӨ�
����s8%J��Q�p�r���'u�`�1���=�a��b����$��JYw����:T�RJ�K��a�]	�����W�	Ͱq�<�l\�%S�Pv�{}| �ś��Y�[�l�E��4s���W1t��е�#��ݻÇ�K޶�n[��7���W�_��:ݩ?��9G�]�t��X�˙	ݐ���hm�mb����s|�Y�(�q�1�*C���tDL����o4z�BL���^v�eq�n�k�i)�5�E�H���J��[[a&��cm Ё�K�J��~�1�|T�#3-�H�h������o�t6����$)KO�7�sn��N��l�Y����bet5����uCc�c�D�����G�2�;�H��QZ�H��&4�~��,:�Q~��ce���+�R[IjUR	�_~��f��,���Pu��r!ל�)Jq���iN��	l�m���QD�Άs���K��~,�E�8��:�Bd3�?�q4�J+]�ՌZN�� Tl,�!n���/��rY������yp�AM��fU�B��9�	�!��#�|����S;�Z՘[�-	�-�{N�͝�V
r[7E�^>�]�Y揹i>�-��8Ss�6|(2�X���.��1G��M˄>� �(	Yo��ѵI��ޚ2G(<���_�K���$פW{6+�A�.@m��<wJˊ��W�)��/��ا�?�+Hx�CbZ�g�h�Q�
'�;h�AS�6������F<�}	�g��W!�[c�v��n8yͫbU�,�>��!�4��� O�{>�Gu�(�b����0�@�+zX�z����kk���H��F�S*O~��[f�ö�����k��%��?��z�����Ǜ����;�=��sQ�ڍ�?b�!��0ǈpD���͢�����̳���������Q��o�����4��ų����������'�ڎMm4!勵����4�+2�f���:����߄�j*��_;�O��B(���c˞ĝ�ō����U�b�i�`
B�H�t$R�{��'ٳu��4Ԋ�CR�d� J̓��6��Uk�d�8����0�~�� ��{n8?q	E	1�7�8��"�`M/L.�I�޿��T!@�h]��A�Ϊ2ݼ �mJ[]���KKnW�0<е�퐝�œwpayr�Rp��.-�7��N��]����K��`�T�!<-edN�q��oM߿<��K��T��˹4C��V��!ޑ���#zfP�F��>2%q��D�@��̣�g<���_��O�tY��*�Wڶ�1��|3�������m�?7�&���~?��̧I5W���<�R�  ��_(�2L���δT����JU��
�d���8��0�R���B�,����i{�҄�, ��c�xL&�d�R*�{�7���H��& *��+1�G�9�rqQN�-Hh~Ľ ��뮢�('Li�,��,��S'�sp��o�W%�� m���cs�\R������8��H����6�����9�����&4j��~�ק���a`����$Y?�W����ă{�^�M�ų�K�h|�~$g�LL!��B�M�JPjPLX�j~w�|���(�~4p�,N���U�wH��/�5�͊!�D��A|��g(���C�A�D!��Mύ�K��k��9� 0�������&��5�������Քl:b�Ϯ���;���{2!�V7�.ۊ���nk��`#�^V�CvAqčg!)��#4r}�������}!5Sy���m��OCH�w�D&������;@943�3|����&oB��p����f���mS4qv�!����A�w]i�P��L9}�X�L�[��3 ��'w������H�cT�@��GAr�(&I_�o[$��B���k�;������¢U-�a����Q%�f�.<�ׄ(�Ƅ�=.�$����$��� ���V��0��vUUK%��"7)g:�G�r�9�7:i#��pD��O� q�87�ϲ�G$s����~ t�W�D�ߨ��*k�n�{;ac�m��܎\��=�M����F_0��u�F��0j�C��y:<�a�\OI
��v2M�ː[vMw(-�MX� ���q��#C��acӚ�t�a�Z�>_����_��sr1�8��&�M�:�Y��4ǓT
�IlV/L��|iF�c�9��J��!G"L6\4 �\K
�&��8fd6��d�3��t �z≳/~xzl K��)�oyV��C�k�N�`���f��+�d��c�(��c���掘b��7�?�.�a6"�S����/U���=������;*�W\��͸����Ki7�>����ݤ7?���ؑ�j[q�-����AK��Nk��N݇VT�8%�P�D]�����v���:��	���n�)��J
�a1j^H�׮�0=�=�.��S M��x�/�Mzr��;�vA�#�\&p`��RFn�:��?�˻���uH!fn�冀�Kq���©�/���I����"�h���V�����"�i�%GeΠ�����|�o���<��=��ǯ��8I$<�i̳�m:N����}K�<hB$�F���4t�v���<&=��͈��~_��v�*З���hp�CB�ύ<b�+��\+��V��2,MmE�<�����tEob*O�n�}>c�����~���x2g�|F@uR�v$��1�ZY����)�)^��9��4�+;I��:��-�����@a�9eUQ<��[�d�(�%d��rd���r<�m�K����w4���ql��
��$��1��&��(r��g�u�P�(��ˠ�J�+�z)�\�)�	�8p$��G ��n�|l���N�vHT��Mׇ��(��.�5�>{��\���4�7�`�5��%�{6!��M9�@���e̴F���z�ڏ�h�����{��9͔���仑J]�(��o��c����*Lk �oTT��'����r]��y�o3��<ʱ�p�mt��r�ڣg�J�1�ᤘ�2nca���C�#���=�֑�I`ۣ�0,
һ��v�%�%�}V��j���JJ�`�(�]#�Ѯ�0��8\�;&a�;��y��\���#��9�r!��g4Ȁ�輁'T3z�y����ĳ��}�'��Nꀮ ���l3|eᅰ�]��f{�)�N�O}x�O�Cd���	�:ͳ�ӭ�q���1j�X}OԾz�wo���NR��>�J��ϥޓ?(�j�3�ݖ�����~W�g&XjnGz�4����V�>��S@E(k�0�mb�D�A��
��)�����o��ʢQ��&識t�и�r�����N� tܽ�Y��D�/��&L+-��fq`�y�Th���M,j�$bSSq����Qg�&������T�-B-��Do�>��o�j�#���|��lت$�8���a۸@2��ށa'���^�	�"z��^����t��@�r�G1���	�*�����>��� ݌ܲK��Wͥ��)t3�֜�qN��O�=�$�Ï>�����!��t
���U��,�$������{�H/�ޤ�s�0ܘ��M��K�R��#��*\��;���s��q���\ 73PO�v�x����ϭ�.j^�������|rK.�{��v�j���۷�핟f�?h$g4�i��2���U���X��T���!�h��9/�Rl
i�"�:�F�8y�SH�EC ���=�b1يڟL��E�<$�N��s'OH��y��zL�[�*��`Z󼶴]&�:��36����h�셙{�w�X�\�I���x����ݱ�)�~8�s�W
�f��:�
�5+�XL�h�n	�;a��������������cqY��+�Y�ݎ��<+��Y��SR�-�@��J�o�f	�A�&�+�G��x�\�����EY9Wv@�F5�CS�h��kTȎaBa0�[��1oH9WH��JZ~e�vHJlg�S�pM=�a�weQ&�kGq щt�BM-��Vd$eb-�-ء����k�T�p*��T�Ƙߔ�\U�_���<�b#=�Y[C�nF�X��J��MSrz1���!��Wl
=���::;�YB6^1g��Aw�ߌ��]eU����Ɇ1+w�px*�\u�㎹W��'>����^s�%HvIQ��������w5�ku�0r��s�	���L[���1� ق��ב,^_�3AD��X�~��暙١!��V�~��c�A�8@M`8��$~�9�B|ri�
��>��$Q�|�>�c��P1��w1��L��b�yڒP���V��C=����So��E�0N0����z�ʅ?::��c4vW��
�	�)�(�ə�j��z
�1�O2����Xb𖎣�7S�9�Y��oc(GC)�6CSX,��/7ܖ�fΖ���a����*K�I���+����a�f��W�����-odɛ�&���[���BvuBn�36obx]l������O�#8����n⦠r�aq/� ��GTr4���^o�X��"�&���wJp@���K0OҲ��J!EڋdPw�`����{�u��ab5������p�k��{�R\\�:����-��Y���P���]�9+ y�{=�M����@�P��b)N�ۛ���+��-{��/��6��S��S����>L�N&�9��xMx&P���|i�N����(�(=����y�ξ��9�qQ�MqR�5J�yק��<(e�:ANC�m��,�u��.:Պw'� ��	䡊�fV���2x�,y�� �8�l��w_ç�X�:���?�]�*b��n���M�r��q�A1�bT�G��ܭ� ]0Ə#�@$���
|� ��"�|T!�>�w�U���y�J�7x��^����4]*�b< ҹ��R��Ƣ'A������.�S��ݟz�Cg��x;�2`%1�@�����)�@�Մ'�b0��PE���jrUv=�X�m�Mԝ8܏�]�pRG����a�u8jJO�?�$8�$ع��
�AE��uF���fʼ<���j"��0jO��*���}PW8��Qw@_�#x���m��!`��D�:0�,쎄V��|�C�G|5�����'���UDѝ��皌	�9���	�~e67�jJ�3�#���(Ӌ�i��o\���Fc0p��C�t�'�.Ff"'pZM"{ "H���5�N�rΊ�[�἖�:�x6�!"���sf��q�[1�Y�:��K���p#&���<猞̎S+��lF�25��5� n����{c�t|�JJ�"�^QǢ~"g��"dx�����va� ��}��aJ�2��
�3�<R�-�3���s~+h`���?"�O�V�<(�����ݒ܏����R�b�,�_������F�/&ba����o�7Ｐ�y�P�@.B�QBo�v�lL�g���荧)B	|�OJ\
עq�^����D������(�!�� .OܫÕ+�� I��)-.*���i�3Ÿ+b�M>��3�"�yڏQ� �+1�[85��^.�8��*'!%�\������[�,��>~�1(N$g=�4�'w��z���Ѭr�_"ZLjH?F$	���+a:�j��b�F:1�ƐϨ���B2�����P���΂Hٗ|D ����Ӊu�b����-��������5Kʳu9�nC5�K��Ƕ��d���#!Q�[�ٕ�c�!e�����DI�Z���oU@T=�Hk3�P�Lu����<��盃W�� ܾ�Fc���S����h5ޘ��nm��#ھ=�=�	��}�t�/���2\���2��>�
Q+�O�kNVe��Jь��P"e��{K�m}m���+hb��_����>90�HG��H�啉�R�5�ܛ��$��h�L7C�;��dQ}��X� |�k���\�c4lC�7�$���c����	�b���D��on�s�+_��4Y:�Z����I�^�p0n`(����q~��I����2�sy���4^2�7��B�i��q� (���,����]š�_<��<)8���i�|��qR�'�'g�NG��E��)����lC�3�����B������ЭQM꩐-;���)��i�;�Z���Q���J�W�&^m�����}��W�������Yn� �!�]�.!�AZ�ټ:J�Y��~':$��Xm/�+�vka�֍N�ľ儙�{�9�xڮ�G`��P��L���"quj��t[=��#��e�>=r4�fگ��d�6)���Fl�R��G������8��t������J�1!%S�\��}�n���Z
�)S�ſ���K���z$z!��<Ba�I^��@�}�OeS�F��Q����E^Б�3��n��4�L�W��Y���B��g�L�4k�2��V�4���e�H���ʘA΄�ű���;�i����G���YD������Ȥ x� �^�!5��#������d�}N�.xIi
T�ݺ-N��&�?J�GU�^����� �ݎq���}��i0�\�UL���Y�;�'��p�b�(��/�"�}m�@_	�9��i�Q�z\�l�!�b͓Ukru��s��.�.�X�Ŏ\�f���>�W�&����=�ϦŤ�`-�y��<�=��yP��-M��p��[ [�R)�b�aPbDh�U���?O:����&�4��X �{�^��g����N�qM:j���;��z���P��u|.ުgZ��֟���_�5�n?�pN`$�ф����r�XU����<�RM�q��B�n�_=��ׅ��٫�q�6u�5�����7��;<�ڽ
�f�bV|x.���Xw]%uV�k!c��f����a�T9T�=��(���R�����#�eRE���
�r�L����޽]$k�D��GG�C��̘�
��?Z54`a�0\x;'�����kA�p�Q����2c+$��7�t�o0��R`��u�ow`k.�q�?�Hέ��2��~]���~��K�������B�*�r*J1U����I3(��~X��Ȓ��>�a=��Lt	�I����BVs!%>?u���x�B��*�o����<c!Q�W�7�I��d��Ȗ
�2�$�<�7Ҡ�l��vV��CH�O�?؅�.gk�h:���3�";~	F-��L.Ģĕ�#aD�E�ZF3yos�@�ňl����J�3)�!�7X]F9}�bUIr��`#�m8.k���Œ)��g��e�[K��+ޱ�
���F��?e֌Ec<��~X틬V�����V!��P�+�C0Gю�D߮�T� P���.�k{�p�����-4�b�4Т
��������)�����[�^~�FAj��D��8�=6w	%2HGݾc>���H�9������x!m�Mej�N��p]?�Xh[C� ,�0h�gHpO�����bn���l���hv��ؖ3W?�e��,{W��c��Kiv�,~�e���k�>�'TGbYtL�$N��T�-ߒM�;E�q��q��XI��<�]�u�x�Qx�܁ňt��.Y��7i�~j�o�0�?�+��2�D�	�Ө���:F"�-��{.,�pS�W1[�U܋�{=��c}&���{u�m8�������1��1�V��y��|�a��j�j��r{M�%f��w�8ɂE���4м��������G�"�X�A��
����4B0��o��9����1�T��l���,9g�n�ȁǥ�|�4E��Q��$HB(�:�m�:�8�0��v�ǝ�^6�6m�Qy�	R����bd0�	����Q��|���x��q��< 1ȭ	w~"�uqKns�VmLT��:ki��*��,%ʋ�aыH�e1l��W&v�%O[��3�O����Z�5K�O�5Jm�z�������F$�iC�*Q�y�\G|(�9�T�h�$9��#�OiQv��#�e��\��8E�ӕ��a�H@m��^R��έ����� ��n07�	�4�*p�
h�z�p_mi��t׵�L���r2����1�rH����e��'��i����Pz�c�4>��r1���V<蒾u�1zs8�j7�O��O+W��~��[��n�/�����fv�C����Ҟ�ݦ�9�GP������Mt�y��g9`U����ӾO }�z6�-������&�.�缡NtM��S�.�������t���"���d9�b��|���(�]���no������� 򖳵j���$�&��l�jA�Ó7&Ȕ���8A��n����M�a�*��QC�����x���&�xv��kn�
���d��m`z(kΩ�{Y)	�'�KŶesyI0�����{E���%Q�x#K�VVVU�Z��dfX/����3M@�S���r��?u��\�v�����r��AȻ}uRm*�17C֯FUz�(K�XO�~zN`qL�	��C=nLs�6xӾ_j(f�{#�pڽ�zo<���Χ�L��%p��;"��/���&(gFf���������T��]5�x~��mU��?����ؽ6	q�	���+bG,�.-(��<I�PqJ�,]T��a��d�:9d��W�r\��I~�n��I�vS�c��X���Z��;�I�*�U�D��V�(��L�.��L���ܓ�u�u�2�iF�Ո�v� �.$�[��d��Ǽg��3��LV�L�ڴ���5��I$SD	����C'�kT��擄1xC����(c��^��yP˩d�ͤ��t�!A��B��_9ߍ����ؑ�vP4��®b�o�0Q6>���$���1�=�L���x�HZ���@���"�h8픒�$����|��ye?�ۨ�Xl��7Dݣd0��<M�6d`���r�n��Z�9I0$jh	y���$���+0���G� ]� E)���{.,p�1UP�������+��?�U�@AI2K��  �S_�3=��;]�K���j��ȅ� 6+�w�0׼N��U��n���-��Y�y[F)g�#���]œ�H��l���t��әGK�QC� "E
'��
V�ƢɁ�/�~�4p��� �B�B�{���$��R��6��2K1�ҕ�G�"�g���u�^�Rb�Bi\o.QS��o�St;�@BԱB���)Q(�P�tb�a�R@���F�H��
�/�w��p��^�|O�xk{S�h0�g!ik��w�v�va���В�6�&�?Qh݋� �
�����u�gڡG��w����ܧ}�C��jy�u���k\�C"��j��B*3Ҝ%�J�����@�?��&�Eg$�[��;3c������>.�
���O��E�X�V�vϤ_�n�ȍ俑sƺc\��Ǔg�O|H<w��P�W���v�i!|8�/l-��v����t�a�p��$�����:I�Zt���)!�J ��?.��[��pP���[)퇆��h�O�,�ι�[��QJ�^' �5���a�`mUo����A�e��L�/�X&������1n�v�N�(�-�b~�M���Hv�.�ѽЋr���~�`�_�n�Tws���(n�������CzF��W∠Vh�!�Pf�e/'D� ����Mf�/=aH��,R�Q,˝�x�O�6�Lh��U�L���B�&t߷��%iWR�͜�㕑l�/!�߉7�^4lj"��͈�����|����^d^��áM�<4-v�$�ؔ�~H�'tG�)�M�Ɗ?C�e��;�v@>I��&�lFi�)ܻܙ�j�:&`xԨ����l�u���E���{����d5F��G��۫t���+<6��vyx�9'�s�W�l7x`"�'d����exS����Է�T���n��.�f+�:��
�ju�KJ���B����Ju,�οb.n�[�^4a�?_�.���=�N^�Gp/av�~�}8�����M!q��.G��oUf����?�=k2�V1�G�]�95�%���a��I�j�s����%A~U�
j$�c��sp�s}υl�� lX������Os�hKY�CZ�ǻؐs�?v��s��1RR�M>�>�|�L[!u��pLI[�ppm.��]��	әV`E2�H-=ƈ�~z"��N�����gSV�G��J��@i|.���x|XR�d=��1F�Q���m��,^-��k4i+ݟ�ˌ绡�c����"l�7[��*ҧ)�ܽC�?M�Y�G��W��*)���(B�)���!�?���z��	������%Ka���˓�F�/�K�	����K��ee��yaH6�Q��s��x㸮�F�F��*-:v���(q��Ӣ���ړ�p�5�f�����AL�B�`�޽ò�T��_��&��,LX�>J&��R��qT>�3���nJ�o�ф�E��9���i�n�j����|��k�eZ�N����;�^����+M����Q!,)�X!�?�����%>:�9��L7{!f��,��s��b��w��H~1
�̪��<�a�R�$������������=!�~��n�NO Ȏ%�3FMn���X�!���V$�%)���>�S���A1j���s��%RHNoi�i{�l�����_��Eζ*�?��IF�����/��n�.���%jL1N�!��q���?�*xE�k/������_��/�q�CO\f<J�8]��q<0��4�3��ྍ�a�݆LƝY�b/3��=2��y��,`!�Q�1.�ķ%�B�
U�����qV�KGN4���ءl��T*Ku5,5n��x!F�N��1[�Y�'�lNiQz_ޕ��n
?��"/%J1L�g�h�(1]*@
�^#��$�S:��B��J�n̷���y! �2@܅I�bw�����(v9�*%C3���Zg�Q�cDBKM��G��r�NŊ��[[\�dx���qf�!mv[�1WAU�̖��{jz�2wo�k㡿�;�1��
�H�и�痺��?~�/�6b�FS��6�Q�3�X�3�}A���Fkڟ<�А/�7tO���m_ZC�^PI���P���a�wP��1�2X��m��"�	����֪'��'T�v���Y����Brn�FaSx�q	�
`$��p�2j۠L�*���ֶ�\3�hI��v�)����d�Qڋ��Ua�o�c�O�$S}�1��vv-���n�#�r�~S�&���M��2�Ǯ;�no�e���&K;�K_?AE���̃!�W|��z�I�U.o�w}����}HZ��)j�
��$��@W��T���*��Z���0�wc�����:��o��v�	+���%$�9Y*Fw�T73p��!R�=��� 3����������I"�R�P<;@(��Ӌ�p>��C˒;Y��}�/..�ƪA$�P�*������D�2n1�9���'����82|
��$�CC����q���j��Vl=� ��J�v��c�V{�0�H7G2uj`����s�ȵ���Ш~�{\�O����0b'iRrX[%�O��9���Qw|D�#&Q�ɫ瘅^�I�~3���T��*\q ��5�N�-
�_�g�j�e����nv�li)21��s���>GJ�B-����\�u�u��±�m�cTq1��������t>%dȈ`m)h��/�A�}@M�J[�<G��,��.}�!du��.Q�$X'���80b
[q�]����ȡ;����\��NGr(�O9�r���I��+����Ec�[jk��o�!0��j�jK�z���iwH���˜�9_'+�M��'�XTc��%\�۟���O�Zt\xڲ(��4ac�Y0`Yg�Kg-ͺdR!@���� �ĥ���W��3J��
x��(�X2�t�]��1�p�.&���S���wr�EՅE�����9���֣NI�Uo���x5�śV�ŕy4��}u�M��2/�G�/�عM�X
�{��"a�UY�>�^�"x���ւ�)Ť��`�����VP��~��w
|7t�[UT���wN�� &� �h4�l��#��Ï욍Di�ֶu��&K�I��3N^P��n��!sV��s�� �fIX �9�q�I�ď^�.�l	J{�������[�����ݓp�G�
]��v�ig'���"H�����J�C!�K� ���&i?׬&H�@������.�Y���wk�|�r{&T�"A2�{�v��jX��`B�c�p�Cr�0k���n8��5����6*��B��[��'����#�~�aR�~K�����_"�3������S����l�p���ܷ�iSG�`��K��%��2���f܈� �]	�Fi���T[Wr��'��D'�p�׵U��L�_�Ə�5���G�tO5.^i�]�X�,���@r�i�@�q:E�ٺG靁����.1N)hV��@�E\x�b��o�85�އA��l�m���	T�m���8�E*k\o%w����a�p'�?�����K:]Ώ�Hb�=����>u��E�����T�l�߇ì�*g�v�A�m��Pu+3�:�n���r&��k�i�8��m�~@1�BWý 0IK�v\M�Wǒ=�����r؁Ej�,�v�F�lW'*�f�˕��e�S�w�s�O��%6�:>ڎjNU�A:��,gԿ����!+�^� �0ĩ�1�/-C�L1�MN#��"� K.���9��h�9F�X��6>��pr���[��Bخv�=~�\�ʲso/�O��\������E���L��p�>�85Z�)-+�wA���u�K�;���ķ|�|1�/��v�,�W��˳(�!"�"0�	Ӓ����FnoB�>A�(j ��ʭ�POd�/��tZa�E C�x�洓jH���l�
j�t7��u&h�E��K+�63��T�� �߫���jMd�X��&j'�X˺�%�����,��G��|(cɺ%8>o:���hr�@κs�3{!�v�x����383{M��ǵ�ȼ����l���˳uE��e��kG�0��U����ȤM-����2T�_������L)ȸdug�������U��L,F4t��|�'u����ʛ�"����d$��p��L�OK�ͨM��8����	�%k	.j�;�A"��YO��j)e*���G+�V��G�e+o5&}f�~��$�o�vZ���XY�!D�f_ ҹ,��t�&�p+��@�
�!E	�a�@J�C7Ю���&�G��Ƕ��-�,��
�L�֧ �.�4��/��ߕ�}���hR�Dh�
�9;�*6zj��M�t��E�G� O�b�U�/ɂ��&I��V��o	��y� ��t�$| ���<��ҽ��)�S:`|�؃��+E���@Oדp�����2���h��\���H��`ҥ���b�:�js�����'���� �ߥ �Û��-�q1���F,¬?�#o��!��$�qq�࿥���D'3��xlRO��D��ە�m��x��
�1�VAj�p�zu���eQњm �\B!�||�]��r��΋�h��h���䵜�M���������ٟ�f�G>B���� |Gj�V�U���~#��;�^Ժ� IY��1t��}�J�&
_�k��*���s��Gc�85�ٍ�Jm��1)cQ�BH2?ڝ����/�AT3��7퀥�ZƘ�(ipF~��U�X�H�O5�7NƊ�r���-/[m�b���ʳ$�ѽA���4&�+<؋i6�. ��"���ZD�����&K`2�d4�:�t���0�C�xσa+i����܆\&�6
�:B����P/ԻH~m��	��\II2s�Z�B�aN^R\^|�9�3ߖ�^�B<�{.q	/�vT�Gg��@\X��R�[H�o�|� �vC�֣��T_l�L���iz�5�������G�a�6���;৩45�K�n����ɵ�d�R�o���C{�F�k��l#�3���Y����4'�Q��8���Tw�T���c*�I�Y6���Zꔧ�P:���t����-l�Eյ�^r�s }��C�1�5SS��ݳ����,���3�(��Iί>
Fk-(�P�&����Bdu<���dO���e�j_8��i�0D<5�_�E��p"��+y�R I��|�-MO�ݹS���ٞ�!ZP����g�h��8P�H�(5$)]?!"���y,)@c����'��	�3RhgL��k�-�g����g�}��ʤ��T��^�x��G	���STH���k$)��4\��] !Y�����>¿�>�#v}(�+_�lȥ��E��u ��׷�K��e�l��OXY�Ԓ����}���J>����O�M��};�v�\d���O��.�E��y�5`���iFN��A���7E3���t|Aƶ�	����C,��]T�Ex��fɫl�љ���0g������+3��H����4�`���=����|��ϯ)k�AV�7��Є"��}��>���U�J=���E����7qW�Ҷ�	����s���~~�슲�K��HZ�dK�D�8�����Tl}tI�`38O�v�Ϫ�F1g�~����ͻտ�K��S�`ކ91d�t�z����H~�W�䪝]p�(�&��ö�Sb	I-��|����5s1�Ɨ�G�J��|ZG��K�h���t��&�q1�������!���Y*K������׎TR��k�����T�4���	���s��[E�.,Z��m^[�`�oHH�z�X��9=��l�f��z�
Cc��1d�_����jt1��n ��o��p�]�!�����־l/�<c�򁪰����l'9���g�1Y�4d��X.)4�'��l�m�	
zGR�u� 'cP�Fp& U���z�,�zc>��o�o'�7�d0."ٲ�-!���w8V�K�������4�C핡��E%%B���,t���7���YQ%/� ��|�t>$G �~ۭC��b����Go��Je�z���>/��LL.��И1� �Xoa��� ����_y���<��VE�6���'�n�_UXR2�eq7ZQ�Y����:�7�h�j���
+JFoN��eU,6|g�ܡ�䉬!|pm�q�Κ+�Cv�����
8,��]���_*�ɵǊ⻏��ѱc�{�jtF#U�;�l&7��o�@X����Ix�~v��!{����=��kf}��o��g@C�nم��p}f����#�+�������2|��X������:x,���zT���]��w/릝�8���'L�O����xFk3�rT����E��F[ ҍ�fa둃qL�r���tg��蕪p�X�Ǩ�@��?GT�����)$g��3�3	���䤯[��q�kgy��V��E�d�����ӧk�S�3~"�������AD)sbo#޿Ƥyh�u�c�98\Xt��� ���5����-��l���R,-T��w׍	����U�F"���'�zE,�o��<w�Iw��;D���5�BD�33/Ԉ�eM �4N�~��z��RZ�,RH���}��:��S�ߵ��	H�dG5�s��9�U�YAC�ܵl.!#d�
V����Ȼ8|�^+���!�D�����g(�Z1���������D�o&�{����{ӎ��Χ<�b�7L�P	^I���ۿE:���SZ ��Uf�ArfeaUNC2���T�����$�[F�1S2�-8��Y�!���dS`~��e�R���$�-�:�c^�T�p� 9�~��:�6�4��Lvh�Ւ�$��	3`��5[*1tC�C'�c�Wd)T`S|�B2��%��G"��}����Sc-J��
�V�[��ΆU/����FKLo�M�~��}�)F�n�W���?��Ί3�;.ˮ�?{�Q����ǣ�
̀�|-mIp���ʏ��	)Z?y���^�6d	���Z�5(q�����tY�3�E&:�c�8x~�B��E/�Γ���Y��,�I�N�X�z��!5ҿ�\ ���K��Yv������^��������H������S�!�N�:�	��0�?]t�2Y��u!����hg[�(e����[��׃�C�X�qz���f#�S��f���(ؼ|��,�j��z� �f��9E��j���+��'�Ty9_d���z��u�E������c�Q~�	��NL�s0��rƎ�ZϜ7���U�\B��c<s�6���N�����ȭ��2~��3�7�6�vX*ԑ1~%��W �X�{%^���[@�@b�G�|e���}G熨�60l-c�@2uʍ�����E�����;�� g��7}"�@��܇�~X�&��!'��\�>����bϣUj�gt�;t���Ѡ��x�B�>��6���!TJ���1_��(Ϗ�ek�Ik���^!�A�!n.gqc���n]'��B}J����넏��9��`XM�o���6j��I����R�4��j���tW�MElr	}Mg����YZ�/˞�q�]�� mI|��^.{�K������� �e��	�s���2Do�h�<���[��<7]y^�ߍ�bĚ�������D��c]^?�*�~4ׯErT�:������e����:4Щ�%j^+$"����]��x� ���9�����|��.0U#��h eTlt�KUg�8��+��(ӹ�,yvoo<�vb �ٰ=w�e�7�2�=]�+�O���;5� ~-o݃�cF��K�g��bE� �;6��d|��C>ߒ�X��{k�H&��<%=�TG���v��$�2��i?D@ә�z��=#wa��{���[�=����k�C����eߔr�i�2���� �?c��f���B�VV%�6�)1�t@=�<`#�Ό�3ƨaؖ�6�)W��A��-��'�=�Ç��+K%q�B�z�1J��_�c�Y�����3���Սi�ߍ;U��#��s��ҐO�-�7�gpO�Y������B-k��RޓńK!g��h���#n�S��0d��)�W���y�B���+���0���e�i�jif�Q9-r�� ʟK�}�|BJ��͛��3��d�����
�h[q��-=:���n���hʓ59ʦ�T0�tX�ng\�Ƞv$�ʀ��l�OI�,7$`��V˺�Q�����3��(��;>�"�@bN��L;�>Ź�ܜ�Ao5B�>���d	�o75h����c@1�kp��hl�<��i�Xm
7˰�>3�u|���V �����"�"y�O.��J<����Eh˾:�rJzW��6�pl�+�A��J��j`�)-x-,j�FNe_֝.[�q�	�%���0��ʐ���y|gA���Gw�44Z�x�]�v�yq�"� �:���p�;���4'�F�ړ����j�`�����(�Y|Ի�e/���,
�4h.5�[�TIC��o[�P�Æw�Y0Q��i���k��l)I��2��G��wT��c�{�*�Q;�q�Oˬ@�W���q�7��̉����(�@
j �vձ�7[�ϜrX}�<4S�(ّ��(P��ZcvA��ҡ
��g�>��ۥ�(�Oį]o�n��Xo}A �<���IC	G�i��� ���!��db6=,ﵭ(�W}[��@�����8��y��:�?4��'>�8�EIE�)_�������pV��g=��0u��\рz����<ҳ�NF^h;C�<+ ,0[��h���[��vF*9͉�Gh�X)R����S��%�'tLw4���e��c�0tGVt�nv��\){LdKP�F�8��7�Ո��zWQ�`D@3ê0���\=F��`���7c�1O8�����z"wJ�����jo�~[��eү�6tP���T7ٌ�1m��!ԓӯa����"���n��G��̀��q>#0���Q�eF� ���� N@��?n��#$��h�v�|������fƴA�B�fXٛ\�QS;b"�^`*�F��}��o��1���P7�i,�;:��fR'��Y�i���fD��p)T���j�DB~H�̮+��5�_Y�wA��iv�Г�Ҍ2�;����_��ƌ�Н��\}������`Lh�:����K p�8#5���l��O7X?������ci\-<@x�����c�>�4��^��\�)���=���9����b��P��{W� ro����ȗ+�h��='l�]�����*�F��t:�w��R�Y=261 Α�k�3y��-'�t����0�eH)��R<o�@��9eQ��A�e���T7wْ�	[?z�4��nj�D�$�PRN��*+6)B����mB�`\O���j�R�ԃ��o����i�� �r�a�J��I�O�@�s�E��f=�+�~�K�tqic����N~B���z�9D���Y�i�l^B�����%9��j�$ﬤ��7U��݊v����3���l�zMY|n��+79�2��S?fa���@�W~"1�GJ���j�6��<wc]v�C|vm���=�$߄%��h�Z���mU����@�,gZ`]uԐ��F��〶��^h���YIL5$sò� �]�|��jl���yJ^Zս����I����)_��
{�^.'05.G�2��@*�� �
�Q��Gev��x��b�<�T���/�R��Dq�g�f>*��@��rL�(�{Dンw�^#%<]�Ohԩ�{,oђ�%هfx�}�γ�
~G �>�I�+�2�S�t��Tx��><��	���b���C�n�1r�N �!��s��F��t��
�E�,(T`AMb�8�{�0�y�i�~h�V7h��,��gx�!��dv��g��REၺ�!�dK��V��l���R~s��t��D�arx��Gt!] �V����~�h�sn�e3����!��֣���$�vrCW�d�I�B�	4H~XfL��$�du?V�n�H��F�L3?ٙ;�۩{xv���]��M��Xϗ^|q����lpp<L!]x�=#QvO�{L��*
d� �pY�^-Y7�{p`�7w�&Q����?��f�3�ޘO8Uعo*�c�$�CXkw�/4p�����?(Vg��"���R ��z{��6��W�r�=�+ͻ�ZF��Mʅ�hK	ծ[DNW@*�.�	,9��8���� �!���������o�zI�9 M��K��`6���%�4��DN̡�m�&<5LD��|��HJ��G7)WD��Q�B��8��{�Jܯ�B)�4�\~�z��~m�b2�#?��f��gu���\�K��<���0�k�%�L<19dx��TM�A�K��Un3��N���P�K���H%�_��F�1�)"�o�/�����C�{"8�z�r�:�.�x�#3Ro�7P�]�W��?*;�<�f'��'_-��q|���ry��@0���.�°ff�5OV�"p�M��������Y�Y�D�~��E�(0}i7#\W�!�[�x������r�����Pp����*���i�(E�Y��\7�i�1L-�a�enp�A;� ��)�-`����q��V)WI�*��{^oJ&�\�;�Ic�=��ւ	J���'a)6�9�,�w�[$|S�����n�9*#�"
�M}�U��	b=����tT.������E�lKF�kG��,���=8�H"��@��&)��_���&3��o'?�Ex�>�n�$�Ҟ lyg@z]��\l[�u��]�U@�\�.�,fl�MM�55�\^�h=�_��!e��\�KF)�{ЄRMx,z*,���(���7�Ŵu-m�8�*��,��<U�eKLke��C���N��E	��ֈ-N�����`�H'O� �Ґ��������
w�	�Yk?��AdF�)x���uEq��P��C��3N4��:��mcL[�\�f��5�s�A�*�#�y`��zV+I����5�ݱ ?�Gg�s���h���_�cX{�lk�c �o�i�Ec�-���g�lx]�:r�J����^4���]4t%�O(���eϳ5b6}�F�d�cF�w@I�x�mji-�l�>�UF����
��>����'�gg�Yw>�U ,��ߞ~���$�8o���
O��1�	eк�{@�b�mRr�V���Yv`���!��U	Z���ex���H6����98����(�RI�� �S�4����Z�G���S%s���|���Q ��x�]�-�`��1c���˚a�/*�ۿC�.��x,��r�����d�a��K	�xQ"\��ޙ��E���چ��Uj��1.F
�~�慦��w�<������0ơn��%姚��,�_D�����Q����X�?�34W,~]' �v���o��L2��k�tK�ܕ�k�d
��I��r�R��n��gi�$!`��<$��K�ҮIƁ�O�Op���t W�A�����(�/K�3�J�X�����v9;Gq�F��F�	�)]����)�<�����Q-�|vk���1qo�0K]���]��!{(e�i`���2��(r��*��#qÉ]��F�����ܗb����.��b���s���&�<E��SJw#���!mXh���r�V�J�&�lSܱ���J{�(:�R��#�ƦO|�1�msu/�^��j���� �.�_N+��$y��D���û䥻�YwX��% 	�QS9�F�����.��(f�U�T	���q���rID������7��M�&�_-B�qQYdr)#f�'M�]=�w�VmY�#�ǚS�Q\�ek��Ϝe���ک�ҩ?�����CH��s��G��[tKK��ҋ��q�)�?����K�v�+�<6��b��ࠁF"{J�7tB!�@h~PC83橇��iV���oV�C����K�p]4B@Ј ؋��������]��3M�g���TO��`�g�亃5��:OVX*��{ZQZ&�%��)�ڤ�H��M�42zf�5}t^�|?��D�s��c�W��v���T�[�b�DC��ޫ����/> J�)+�GԦSKBN��:��,8� l��3@"$�P�)a�\��Y��M��a���`t!�s��d���$,\_�O]9�H7�L=� �ahJ��$W[/��x����<kCΙ�ǛRٛO!{gY*xC�+n�fFǳ���)z\PQ��V�s/S�0; ^�Q@6�P��O��1F`����"�S^�%�ҫ0~"�!d�*�q�֕م��qy֖����n�t�l��ڸ�b��_1�@ƭ��X��<��sf�Y���ˑB�e%r�!��F����:k���?�[�m.=��[�k3��E���0��B�Y�:�2Nr5���ŝU��R�"��U������p~:�'����~��O`�s0��B�E���Xo�X׍���3sW�ƈLNp��������T����D���Z�F�>�U��k�I��]LN,���
�Z�h2+ �ur�gF�f�Ma��-x��NTh�_�H$�`>o��º�����Sje�3`���m3�:������S�ª���̩���sґC��w��{%4�BIŌ)Hb���	��_bf���(2HH��/� ���<Y瞪���_�)�����D6䃣<�AD����kr2+uu&��R(*1 �����ze���|ح��u�' ��Xf.����:���%F;t��� ��Süt�b���(���ʼh�۰�J	ۡ�G��V��؏�Յ�-��g�� �X��ZE�o��o�,uh���'��M���뀁�%���i����;����Q�.�۸²�h��2E��#ʎ�A:��X�7�U?0/I��HsC�vBe�R�d{iIt�m����5�7��C g�#T�H�B	��͹��e���Mm����� �}���q�G.�v�+lT�#��"���+t.��B�q�j/%�@xą]P$�[ő���ݦjdĄ�?�\cS��|UUA�S�ۯيpI`�Ɍ�D�\����C��&J`��P=�/yxem�D�4K�?�j.#6��o�J�XaeIo�H,*R�rN�������$��F�.EY��܊`����d�M�&F��>ә@o圻DeU#��2�6N�����RW/tj.]�f���aGG�+�DN_�ua�d��ݰ�4T*���j1�����H P����RBEp%q<��r��N��"� �c��5�y�&�_vn�2k���8q5P��.C���\���E��Lሽ�1�V!���q�3�AB@?==��G��yU�#b�CtR�݅�	�R3���r��aΨsr^#�S����{/���?Έ�9�6������7��(K�Q�S��E6/��m�`�~���zx����	 N�!��ML:L�py�3����3������?<�E!z��d�8nֵ�\
�V��LEܛ�J�	���cu���yJ@s)��QL�b\���AR~N"��M��Z3L�C��6^��5�m�V�x���1���.A�&�l(�������i�+�a�,�O�Ů�#c?%V����Xu�.����K˔��*z�\R|M�р��Y��V���K�i��?M��3��-jwF�@:������X����=��Sl{��%��>�}Q�E
�r,�*#�S�l�I?D)ꏞG��sD�� �3\j��;����o��ǣ�A| g��1p��#:�a���⋷�BOh�A�\n{�p���fĭ�U���qjk�1f��޳�����(�)�i�R�%�?7�q�D�����o� 0eh��+��i��Y&x�����_ߍ�<�Y�9���p�?����0O��O�8T��Kpv4H����y{ ��r��.���}T�َ���b������)�=9h4QėD�;�<�4��79S7�d�:�����:��=5�* (��4ʘ�|�m�����rSA������sQ�V��!͡L�*�dQȅ �ۚR����Ʒ��>`/�R�!#k�q�M�%�&r-���i�n�!\7lBhyw¶��J���`�aS1��V���Ju�1E�:0u��L#�Dđ�7>�ک%y�Le��������?�fi� SA��P��<���f�n�D=K+�u�ʂO��0�ǧ����s�
����\�@b?4���K�S��
0��;�R��Zh�O�8���H�ŉx� ��p>�+t�An2jbQ���TqWdV`�y�IԈ颾ʴ)��4�'���I�D�a�F�?������%D��DP���Pp�Gd�إ@<^|��Մ�Ϯ����N�����S��d�K���Ջ_H?{����z��6=jOOT�F�4$~t��H�^b+i�_�r�≇ �ͭ�E7q���?4&1I(�I�����ȷ���s��ѭ }��2��G؟�F�����t����Hӹ����\������]40��Y�=�W|P�r@�7�>�M�q���U}5����qK|ޱŹ,N֑�m�'u��HцpҐ�R���7"iOKD� hۯ}���sa#�`��S�J�gA�д����ơFI��Ȧ���\�D)�ʍ�����x�z|4�]á�Њ�%�7�Q� _�S�"V��j	LbWB��LSN�;?Gτ�ū�tՏ��0�}9�T�}�E|�	��qCg�~;��m����Zf¾�_E�;	�P���H?�o�%�>K�(�R�ֺ_�J
PM�P�p@�hs� *�����w����66��H8u���rJ������1�c����u6�<��?A���k!���(���	ܬ�g��T"���q`M��6��Z�x���u��iZ�o[:�L���㬜���������kGZN��8�=��v�z�S����8>C�V-��e��B�-E.�^ԄL��a]wS<�b���Q�J�0^25E�!`Jj����?eqM�N�g��������;\�"#�'n��7fBۃEJ�{b����R-K{��DW�l9�� ��^�$·F�>]J&&�2ݾ� e��79���^= cM!dcT�_Q�N)����X�E�|��.�a�v�&؟����-x?�٥Ze�N���h��:|��\�{���4'd;�m���$��(,�Ī�#����1���+��|��3.���m\��_��d���z�<�v�BoO�
��~&8xw?fԴ�z"�8�)2��࿅#}~E���-F���9�yise��)o����_��)r�2|���F�c�V�N��e0m��)}đ�6��:�B�����q�^��:�
E��%j���J��;��k��	����/Hskn���(�>u~1��`�-o�p����pk�t7��9��¡)���I.��cf��[�\�jy�Y���<q��
|kk�j�Hω��8��.�1�r�X�_.�M�ٍ�����B_�^ނ	�M��K4����v�틥'"w5���~�� C��;�����@���A�\lc��r�kAH~�_P�}�ᄨy���S\;F�k�� ��.w�����۩��ZL��*��@W#��؜�6���c��_�L�~�r]'�A�w8Qs�B�)�r�?�誴Ȳ���Y��9y�7�]^bF�&��7z@C&�I���ṫw���h�A���:�*8�W�ט=�d�e%%DdRU>W}�ʨ���s��Ԯ!��5'Bj��]A�=c����y�j��9�i�,&��2��pH�84=<��J\�h6fr�>�N*�ΠtUb8��7&7A�Rgϯ�.q�uJ��ZZ�8	65�`�7F�_��}
>�� !���ȫ��9�SO��꒪s���GqZ���o>;"6+n�G�Z��	z)h9��6w�|Ѐ��{ҙ��\���P�`C�`���8���2�kA �C��Hw���v�=���Y�) �6�*0F����Mm$��jJ��:�Or��#ܨ�1��߶�8􊵋i�	=����T���g��r�Ы���e�@�Q�mw�T��p�m�>��>�6�+H����0#]�g�uC���7M�47����<�j�T�9Ё�őa�T+$蓨����p�mD�#'�K//�m�y��Z�G��6H?�z;�����{��p ���}� �uO�0D鉮���k��1�g������0D�>^K,����v�U^P���6p%��ut%�xT@KdY,*-�ʱf\;�+��P�p-U�CoF�FK@��|z���ƒ���ŋ�x �H:�m�$_%��~(����
��6	�1^L�"�(�w^C�2�y�VX�k�����f7de[˖��Wa��7zz��1�4AJ��=b����xʼ�����ӵv[���_�+���������������K:am\�Va6��Yz�#�T8[���jq��]s�r�� �z߈r����eD\��<�������^78,�ガ�R�v�f�	}g��E}�.�������_����L�KH���� �-�._��a�<�P��U�m����hI�O�\&��s�O�q���С;u1�㊃D&K�����ۨ�J����F:Җ^a���_
d��*���]�{穐(֒�1��Low�c���������ru�~T�������0^]�DR�824R�Y�>�}`C]�PO8P��p��BDk��ڭ���n��M��{�16Y8��O!�۸�<�J��EL�������g@���˲0׼`l�T=�e#|��"{@��
Rj�K�FP�6{���,���ekb��
���_gV�y�S�e�9"�H�4p���*WSy"�27���}�Йk��#��ps�x��?5uj�Rr�������d!���~�[�7�T�f���������ǐ0�ی���6�^����j�At?xJ/8��Ty�?�����L0 � Xe��U�Y����I�,���|]���ĩ�o�ꧏ*`�[��t�1��ڦ��W���H�E�/k�����!�� �`2#�f���J�=�]�4��/����mJ��~�?�+|��T��i�m�"7��"�+�y��@W.�%�գ6���94l��Lc�oF(��V¥����(��r�2�1����O~HH��;.���eG	����(�Srrjd�=����nfq��="g��	���!f+WG�����.T�w%��+%����n���@��C�Y�rt��.��':�gl��[)�*#g�Rtc�]�wc�/)��qB��gk�r�/W9
��&�]�����V��Gy�����y�lB�lk�o��
��灾('v"�1�j�j'�3��ύ����5+���3QI�؄^o�F��J�|�ٛw|����h=���ʸ�6���u�� �_K�Dd�� ����~Y��ؒl�r��T���+�f��=p��t��1x�_�Z:�l�'?�O����t[+��ٺ����E'�	]�hSc_�&i�����A��X���D�: O��n��<�.�k�_،cLLO�^����E��ވ���נB)���f8au��h���ī���E.Ejq#�o	�do���&��������Έ�g��9����T��S�)�X���X�����2�I�s5h�NV_���vd�1V�K����aB9lʇ^�HS)G�J}3_혒ӑg6[e�,���-��N��h��V�B�5�3����|���U�g�־	pέ4%Z�c����~���/x��|�wς������)�$� ���Ī�!O��⡽$LZ�5�VM����q�XsQ����5j{󴔃xˍY�9�����#�5=�N��!B�*fy+��i�F�8��2�6�6w�cFȹq��ٽzVEN��
}�����ԕ�����q���e�ߗ�V8�4<��5ד���w�������Y^7q�6e�朸�!Z9pf���,����U��;�C���0�k������b��ì�k��h6j�Q��."���;mk��Ο�l�Y����%�.�9�z�I�a(6k�^/����C�ӛ�q͋F�+u�3���]�vJ|�H�Qi,S�۠;l��\c@ɽ0��*K%"�x{1E�^:��>Rq2��ձ��j�s�'mhX��h]Q������p�v�&.v40imR@d�Q)yLQ�4�"����}�G5IQ������Q���ێiߤń�4��C\r��=���#�?�x������0XL��决�,�@i�!_�'n���:(}���7�6ӛ�<��E����Y�esN��dB�]���:��@d����n7%��qb��@�h�8�˹���Ɍ+q�u�6�D�;�xzw���֘B����ٰ�~+���O���dWx�v�8�(���>����t��x��3��Pt�}���P�b�Ť_�fpJM�����R�7 iA�~��rU�/�>@lH$UaN�zzy� U��g�l����zj##�Y ��<<3�]�4��п�����DG1m9��i�/��m(����c�������$4�@bC �{:u��M�㦭�rs�:�!�j��� F��ɫ�^�+����}�@=����ٸ�h"�9U�r��J"�k�L?�	'�F1k�M�3˵�QvN��T�����O���kN�/�j���u&ua6�h�N�FL}�1�]����VV�[�
����r�7�#խ�0Y_���Z�~>It��)�Z�M$V-��H
?�:	��\F���E&`�����="�@r���2�=k]}�-/k��җ�N֬-G�J;A���r�̞BqW��?��ve�xF�W�����7�%���a�7R��t|M�F��y]S�5x��1�hS��5ڒ�b�P)���3��`��Ǥ֥���(�+j|�y��J�mJE�iєo�e�P�C����;etH��ԭA��'���ټ^5R+�i�[�t�{��}Ƞ1���e�I�x5��J����$�GUgz�P�z�4��������S��y�,»��|a��W��v�"���0��g��� ��Џ"�?��:E
��~��B�6G|0�D���e; h���C��]؈BT*n=M�
�`��%�Ѷ���:<�V�bh(A*m0n�#�v;*��������f6�:\ץy}T��ȩ��Q?
��4��Q�R'R��� D/��09��k��v��*��S~l�l�|�~р2�Ì޷�"��R���p̚V;L�[������᧱e5pZ��g)�`*���^�����8�4���zB'�\���!
��J�1W��'��f'������$�-�kI������uo�Ͽr�Ǌ����~o�t�d�s|vWRo��a�-����}�v�]�<E	P��΋����e�Jۤ"�wX�C���U)��� �R�d�+.�[FV�3�0������dd������dӹlF�"T�HH��U�ּ���4q���_?#�W��ш3��h��`ß���N���g����M�{'3��Pa�^��?�Cmc������r��/�3K/VX2�%/>�d_�0����cү��xE�Ώ���T�g[#rl}��=��Jq���5>=�ٞ�{ћ�� ��p-]b8��r��� �k8
������%Q����V%��R/�������^Y}��^7o<���4�
��ƅ�%�	,�6���]ân՟A����}]o	{�a�����]���?��}{ļ����V��Tzj/�}G7��!�)*t�J�t��dզo�����lG��]kW�ҋ�PRG�ZO-� ���c^~����ܶ4�$�gv���]��Rg�Vf���{�z<H�2�+��L���N�Ҁp�X�Q��09y 	�g�u؂ɞ��1i�QG�g%y��5Ǻ�Lg^�1
:
����Zv+����O�6��G��+q��/w��v���*d�	�'GN)]�i��&вL��f�M�=[�j:&�t�Ĺ$�0��X���@5-2�`�
����K]uG|��;V���rM��){����$��?����}_��*q�ܛ�yL�l�GM<�0�b�}�f9R �o���6Q}����5�5x9��
z��|jb֏0�����
֖���n��`
�����6�\VcK���fv�E�)�R'���H�YH��]#7�l��O��/���U��^-�p���kdr�b�\�����))OJ����ႈ.<��wjǌ��V;���^E�]3x ���q��#^67�K�l�=.^M�6OV,��
z�mt�0��P�Lp�TH�>�%��S"�]3�?�7Ԑ񓴩��q	��N��H9�7"ea�u�LA�Rea���W�ےU>�;Q��)*n�zs�*v;�����x=9������!�6=����GT�1�up6�	�#����d1x��H�9{������n��Ϣ2#�wws��� `�;�Ŷ�.���� Σ����<F�,��Ew�[�4qq�Rx}�>����Gi�T+��RS�ܴ��L̊]�֐:����x��W�w�}�~�� *2�}I�0�zJqkX=z,�=��1<�3���;���� ��L�c���WUi&D�&<@X�AT�]Q�|�"�y�e�$Lk?�����CTR{�'�7H�TX�{�&�������n�y��Y�� �~=����74���)��؎ �k�:B�l;�԰g�03Z��Y\7�5Űh�AOw@����Iuz^� ��r���R}!j� e�+q�DwWs�CZ�Ê�)O�s�.���-,��($�H�=nAڅ���h�B�<M�S
⇈8]��T�u��?|�E���S�����q� ����l�V�ݖ������������݊��.~.C�G�*�s~w������]���^�����4�Q������jX������)X8���0~>��ܹ�:�|�o	�Iz�0a�~on�hڐG�A���,�#b���\HZ��I��!ᇎ�SL�gF�̆�^�q�^�+7�Ô7҅�[t7\2�Tq���7�&���$��.8gy�{�]��s٧�M+�ˢ��4���3�~?�h�;:Mng�Ŭ=��;t�	�?���RC�����u�0P=�HH����$HjZ�J^_Ƀ�~�G�={����q^?�W���˿���P����l\��tTV�j���iN����N��o�G���N�h�&�ek]x��]t��<����A�rJ�0�xQ_��!놝���J��q�#���:��ү�K�^Nj�b�6���eu�e��=a��$\�ҽ��78R^�ǩR�nS.Gڶ%�Z,i �0�>�GE�W{&�L�-�f�h�['�(�˜*qLSꘖ�����rx�����m2ɘ���ӭ�	�%��m��Y�o!U0vo0��6wb����Y�r`<�%қ�蕮��f��M#�w^܎�3�
!A\�����G�
��x{�<˲X�R����a3 �_����[�v\e���9����?�S�`�Z�cF���3q�F�cݍȲ��>�)2�QS�0��t�ؠ��t������f�2}޾�V��x����2��N�W���z��aB�7�*5ؠ؝��y�yU_:���X�ؾ`�f��a6���Q��Ⱥ�}U>@=�zj���f��݆�V���њ�Y��.��E��,t�T���'<�*{�.�I>a\I�H2NO���:Y�գ"'fU�Ї�U+�{���%��%�?bR�%E�3�fV�<��[V3����.� �������p��kqU-��v���0�rg��|'�1��F9i��(O�^� �%%0�]Z���;�ʘ��Ĉ��M��m�
	_0@��e�.}ng��b#�?�hIP��c$�N�ϸ�*�L����I��u�0�$?|
եFhVvCy������6�Gغ>�Ս��N����~&�LH1̫�̇BX{��Ԋ���1��_�}��{��4\��7I����Ʒ:�=\]�,O�%f}�<̚*�>[A�Б�g��
җ��7���3��z�҃�Qy�a L���a�+5��u����������⪻pH
��I3��8��(��BJ��E�~;��X�c����zG(�2�lgM�)7�$���qcf�,�⥩��X� G�5R��;5I���J��t���bdTh�l2�~�A��p�OIl�.�LUX�ji�[_[�܂���m�kpk�OtUBK)�*d��S�qU�����f7�w�@�g�C$X�AOc�NB�!y���,g� ��8�_�"�ο�+�� :�Jp[���qkj5�X��T�oyzs��}�6�-�@�0��<�TÅ3:v�N�b�����\Bt��� �e2�Do�b\{����{{�,�/��fм$�<����b��c_�h��64�F�����~\/�ہȝ��E�N�� �8���h/����QDma��8%:�����F`p2����q�ی5�'����3�~U�j%���٧�6�[��+��@y�`WsMڒ���Uxt�X�<.���*8K��F3�6r�?!c�d�Q;e�8'��*�y1���e`�2�ɕ^)�Ϩ�o>s#��O1,�)u��$\r"�g.QT+˚J�Ύz7�~�
&֕&���^�:��yxIk%
׬_����HZϗ%q��(�x��ޣ!�ӓs�ꗛ��9�	%��A�;Hp����s�>\��A��:{�6ǣ'q�6��g���EtrG��	Uh���둽��7Ht@jIfl@HwUƺ���O1��WX�d�o(����L��]�זF��K�.vʋ�'�R��7h����g)|NU�u���V�d:6\Q�I_����~[B̊æ��֎��v���4@���X�`��K!�u!��d�c���
-��Ȥb@β�$�Z?h�Q.�;���,���$7΋�sS���f_T���h��d�(|�s9]�K�TrmUG�T'�&E�`���8٦����ƨ��:6�BR̚ӕ��,�s{�ӇH:��(\�/���ƀ�Y��I�5,�Vm���4\{��j���
t}�j-�~�	أ�@�w��o��8��~��_��baY�+��>�'��dU;���-�x���[2�wBI����+ y&��I ���I xd�4$::�EPG�����d�]`S��Y�J��9�7}S��{�~����S��)q�+�>�_�#uʈ�';�؈��n��
I���k7	ӥ�D�+ � ö}��D�ǎ� �ҶLO+�\?��fF�r�2���8��XȊ�����2�I�f���۰���FI0Z������l	��k8=����L8ͥC�O�}(����]_Tv��' L|wX��*��37���垪�BYS�����C���j
&�w�fl'H���娎`(��r0�OS���97���z�V|,n��o`�*Sv�F,�BT�֧�J;��={�(e�3��[���ʅ�l^���~���&>�	�2 Y��!#ne�%:)��s�Ꞃ�!��+TF��ڦv�x��{��w�]�2��03'�ʘ���]>20�ʒ�b�N����n����j1�h�}�.Z�/8F9��y^�/�@L�A�Ĉ8�0
��1f"Ұ��f��V�6m��u�]Ji_�<�5��rYtLe%p�Od��ߍ!>]nbϡ2��
���I�&��%G3<,2lC��E��'��o����?A'�Z��Ř`��� $�oI�5��+���[:[�uR\�\ء� � >����.M�R�u��Ģ�H�ƹ��;Gɍ�ı�l����Dьj��q�onz=D,L?:U�t���F�9SP�\��?��t�9�Zʻ�M�^��QV�^��*������g	o�<՜���~`�W���?����K�7�p���A.~?@ԴR��q=^�����nr�Vs#c.2ޑɶQ�h�eC�Df#`�*r�gm�b�=9]�t�Ͽ��c�����CM�SJ��4��A�9��B���a�w[����n�46�Y�%C6_d�]��
��bU�?ːb�%7��غp��hM��,+���D�O���QP�]w�Ϩ$�\F�y z��䗊Ӹ~�0]�'����WJ�!9C���Q��;+n�U�����]�E�	�+x��`�e�՘� �_чR��Ww[m�0�:�Y�/)����l�1�W
�@��J��I	7��՟�c��s��}}&���x��D��W��]
�$���3���q"7x�E��������w�&Ck���
�I�#p���B^!��,���v�UGٰ}GX��7���̯��k%q��Ћ��hg ���}�nAW��\�x����z��"P�
�����ݿ5^J�i����� ��(�,/�%�\8Q#����FxOqhC̠��1i�������b�*#	s)�d ����G�PQr �(] g�{���lt�WV����R�	���h/6P��ц����T�iJ��MjV��H`�����A�������b=��^U���+��X����V�B��v�<T�p���j��85w�6������Uږǻ����fE���u�]��3�AܑL�I�H�ha�v�ɂ�IO�Jf��t�����/P��SAET:P�]%z�,Q�k P��Z�EDf}������b����8�je����L�&ߣ8m���ڊ��q����:R��F̠'ٯ��P��U�U�N�("�a�JY/ƙ}���"�qa$�Zt$�>k�7�6VdVo���'Fd}\�� y1�S5�Z���x1��k�#i%��'������>ߨ$M�|ON�f��g8��h�FKk�H����G��ϒ�0o��!��:.���j	��	���6k/m��������A�u1�J��v�+��?������A��c�;bLSmS��o;�5O����F �Rϒ��H2P��;T2��[�'��2?~Aw|�Ug�������`E}�B�_0'��^��t���9�k[d��=x���k|�ߕ,Ի�]]�F_�,C[8���c�J�K�C�)tBh<��S��m3�B|���Day㋸Z?���H<�~O�iy�ͻȄ���z������|�-�64��ͷT���I�*�]i��	J$Z��w�����#|�&x��d��b�\� se&簠�PGYzA� ��ȥW�������8b���o�OD�5,�'�~���z���U�o��/�?Eda�h(YtO%K?��Ekן�\�g��r�&rI�cu�����,���ٰ��&ލ�~���_�.pWC�_��7��}w�=xS��K��	�-=���=BH��I�}�~=��0B�Ho����Sd��B�?Fk�V�li�za�ҰC}���߰q���|_����vL.�.��T�#�����uA�)1;��塴��Է9�����#�	�c�x�o
qA�]�>Kq-6��{���������,���-�M�'u�k`����f]m�#���42Q�J8hg�(�`��T䓆��q�ʍ�o]cG�VW�J9>k\I1����*�h��	������D��5P��LM�tt<���L:��&��d|�c�(g��ǩ;
��*:�  a�.(ki���re
��62gnI�C�U�==Ѫ��{'i�v@���vL^st�2�۳���Q'c/�Gs�kCܸ��Ʊw4�vM!߷2��h�& &nFi�\k��Rzc�2.����*]��%Y�ll��o���÷�:�A�5=y�@^�������E˘��[z�>-Z�m|�mPA�5��c�۸c��+T����s΁�x*4��M
���nű���s�HpEB�Db�'|< j����/G��U�^=�T���tK�_�T��`��@��s]�"�֐)Y}.��o䜴nNb'��I�M^���A/���^�~�Ƞ�ۏ�����1a-y�hQ?aV�i�B�	��� L��V��~�-W�N�"Z&���yXK/i</2�ܪM eK1�7�}�R/d1���VO��x�P��e�0P����6��c٘�f���X hVG&xnF�fo|cߎnw�[gZK�zi1��_.u�����z�P�*i��*�f��^(�M3;S'�H���p�|n*B�3�u0���w
=&�}_i�Uav�k��\ �gFs&�'��z9����+m�e0�j��7����v�;�~�b���}E|9K��m�ߑQİ�Y�/����
�z\�B��ۢC�9��s����6�i����l!0�ޓ��]J��f�1lFu���D���w-N�ƣx�ֱw��ω��H�������lVm�K����]���rߤwtjf�l��L<Ӂ� 响l?�I�>%��((�~�m_�x���̉qq�A� �Q��.�\{�Q�������(�Ŵ��'������K�Udu�cu��tݹ��&`�[!U�ĵV��+0'�L}�.��3������RJ� O���`�d�p �H�����B��ƺH��aPA�����3YK�� ��\�w���쟒	�N�п�����
Mdp�',H����a�R:0�q��r��%�<��Sh�����Sy�ߘd��ˑ�^�?f�V_R9���Y�7i ҁ���EF%�_ܰ�ǺPdW��K�u�7��@�[�Ԟ�a��-9���Kr�Ou�\��)��As~1~�Q��k���ы��3����}�I������C�%�-��`���^d1olZU��h�X�ذ>zq�(�D�6������ȔƇ��ᨤ��o�퇄�=H*�.]_�!�,&\�����@��p�(�k�:N��#���[q�8į����G��~�ɱ�Os\��&<O�{�'����v]��6Y��UXpkr	��3}r�ʈoR^���C�O΂�պ<{i��XX���8E!�2P���DѠ濁V9b)����'9}T4�sL�&�9��@�(�� �E���k��[��#�/t��	.��\~��?y�7CO0I��\���uWS�ZKp���x��i?��G�,�|�Ҙ[�~����'���(����r��i����F
��&���D7��*�po��9و�GO���u%�1j�͏�F�"am��to*���\���=� ��Fj�h�P�l��ѩ�7:����[|�k�i�L �z�[$mgnHӻ��bm�(����r�?��x�P>�[��b9����˱�c�a.�.�U�s�|�kcg���v��7ȱ��:m2�R�,��ь��0]p�|heԸa�Z���i��������5�+\n��pX��O�g������%;����@�����2uE9�5�?^n�="�c���ԈS�DPq]^"gDd"��z��Ӌ��!�қ@�7O�	)e=ů�d�)���.Ю�N0h�����V�Bi	�MϣM&�7E����M=��Y�{b�z����PQ��f@>/0BrO/$��3H��#��ˠ��Y��>�����@�ESw#�A}�~(U�ۦ?X��L�d�|hIݎ��cu[����1ˌg����H5N�J����Tt������hK<w��a�ݓ�e�7�۪O`��%g�[����C�&[��(��6Q���H���Ξ�2y>����v�20K}\�,G�I����lN����e-ma��. ��ߪm`~�����#�����ty�]��p�?�X&U�HA�+�=k
[e|�L���V�\�WUf#���@����E�1�ʶ﷧�+l�\0�`�H��E�)�	�JVHG�et�ū��lz�
�3�@���ɿ�(tP���t��8|V�oM��~�T�cbր;�xv̦Ll�ך
8"��4f��N����	m�)�qI0���������Qc�FJ��\�u�	­�sy��c(zs�A:g9���P�Ƌ J�Ѐ^T7�o���\�w���R��IaTsٔr()�e��k&�į�4���?Gg%XI<��-�p� �Zb/�$��&����U�-����E�	/�G�6�+E՟��'0J s-���ik.��U��A�9��_>���=�|����Ũ�eG���Ce���]X%E��ԚYK��e�d�f1rE���N�,LVG����7o<�2�:��9)��w������W`��C�s���!��R�aVI(���L��p���j��z���?��h&̐f&v�2�2��B�j�;W
�P�/������ x~+�y�d	������{�a�Z�iOd� �4��V1��X����N���j"�r�]�/�F��z�أ`�Y�{����E� ʬ��qit�W��� i��WX�	ӵ�g+p�	�i�v�n�4�p�24i0,8]�"V>�u��'N�}�搌N���H��j��+Nw�C�����8ʂ�Y���<���H�eۈ����6���e0~�~ߧ�<���j�P�Q�k[y���P,{��4jh�� ��Հ���Yw8��A�X՞��)w�c�U�9�5�T�6a-5!��n1��棶�f���2�t�G�D���$MV}�S��+{�݆�+um6v(�d"���e�Y%-&� 򡶫�(���d�#�
6W����W@u!9w�
���Xq�?�,�&���J:��+��U�����hւ�Z�J�'T������i`�M�l����6}Ɵ�X�
����b��F������F��;)�Qh��#�,�rI6K]oXcR�sdS	a��^�������0�4׵s�h�ٮ�B�a�|��ۖ4�T�Ȇ���h¸�����
DgӞ\1���#-����6df��Zmv�z�I�o.�zK�Eomd�"�箿PK��x�-P٣��.�=�i�JR@"�j�z0�w�qw������P����\�w>!����_h��=�[͞��d��-�T���z���)=�];���}�D@L��Hy�PhY��;rd�8��y[�@�Z�>YKk�����V��*�M|\ $��.i^z�=~
�k�l�A24צ�����K�p:�Dh&B(S
�:L�	El���=�f?r�
�:�aj��j�����U̪(����2�GԉF��z��ۿ�݆,_��c�|z�LE�d��ҨO1a�v�MS��7Kg�%��O��"�cc�8��n�����F���T���:�Lw2���a���^D��`�C*�v��?*��H}�Y�ۦ���y�?�W��� wBi{���
�:y������k�Th��Q���� ���ؽ�ũ$�d ���H���fI�Q-�?aՌא�RO�w���C��ͬ�L��t%`��+KY'�FUE�F/���I��}f�D� L�~<}0���h�z���
$_��B��\�}�j�?�L�ahQ����j��,q#�v��d��,Ó36�l�"����t�۔��}��S,?A�	�n��p��,��b�r��:¤R�t���H,s��<����T9,	+q���	I�ji|�Q�I/ci����wN����G�v:#�)�#U�RVt���S�jY�t8;��밑[�@�"ҽƅn}����8s ���|FM3��U�<��m�J�<`�nE*7Ǐ�0`4GFx� �n/
QHí�&�d�Yml�)�{�����������3���4/J�v���-S���_�"��i����7����h|��?=�|xE߅ôC2�JG��������>Ɯj/D��@zzP�<E}��^h?�)Bÿ�rzhi���IѧZ��=/�D2�ZY[?ح�a<��m��wU��Q��f��b�īEw?My�ˡ�U������~���A���u�-�9+˟�t���d���6�i�k�)}m졨iѳ��͏j ��4{��|����/p(%C-��&b�|�Y>\1�I����R��T�i��3�P=�7ĦcՂ�E�e��f�Ԁ۸��6�%Q���*_"�5f�aY����0�'t�@"����*,W�j[Y�e�ă9,=asltt�-�^�J��tt`<~p\a���ع���J�	0m���Jb�};���;�H�pb�0:�z"�`��ʍ���p,����l�#�X|8}�K�Qzr�,Ωɣ���
�u�]K~�g��$�@��G� ���Q%̓zAUAQK����c�F(ӖM��E�5t�[
�d�[�1�A��0܎���Q�n��E-5���N��8kN�.��o�a�X I�[+ّ�H�v�.�y
�j��1(��o�(QH;d����F]��a��'�)�b6�&�8��D�ۖ��	���t�-�3���y*��丳P���i
,��!��쏪V�	�V�c�������@�Ӝ�� ���WNɔ���<�����& 7r�����3�����|��:d�|Ƅ�c��1�+��?)�B�X!N�f����$Q�n���bƑ�'��o&�*c��H�K�ڇ���@�h���(�{�����>��%�z9����G:�Q0�)u�i� ����^rM�=��
��_2Z㔱q�~%p���
��M�;6kvO,����n�B�P�FiC�ψ�G��J��^��
b���n2�X��E��7ecH+9���}�"x�@��	���Z���اu�'j0��2i���Bq�U�bۗ�+�xh����Q�m��aw�����I@%aV�{���� bm�ە�Lq��GaʯLO��CZ��G�H�$L3���X�HV(�S7�F����Eh�&�j���r����Moٙ.��:��_��SV(k�8���i���`Ĝ���@���`9�)�������dij��a�,�Tp|}fu��S_<x����&�$ z��7��S�i����vS��}h��Y��R�5�B'Õ�^�s%"J��l��bsXp�]������FI/c^[rC��Kwrx+�>�S���ݤ����y
�]½���������:10�9�t�GF�^]�ȑMa�쀈�g�w讘�^�M�m��͉9!^~pp4�["�%�C|m1%���Ϸ]p�ؓQ��舧~�7��o&ى���5��-ݨ\9��փȘ▆���P� ����,�!BW%4
1�'�P��R�m�~ҙa�/�"�+�qM�r�8i4u#�Irc�d[Fj��z+�`)�jƂʫ�G.��'���S�����H�R�C�@��İ��͈���-`�d��r(��Yp,CH{8ݼ����^�����g�3Q�]�R��l(� ����U�;����>̃���oŪR��.��,�!K�λ�݊�gq>ޗi�[
h��#�h;�*Y>,��,`N�4�2%�զ��6	�_��-� i*}j��j�ۜ��)�Mx	<=y�����J��7h�'!�z�,ȉ�����z7��Uj�s�0��Q���0�Z�G}^����̵ $p}�F����	�E���U����"%�C.)�2����$4'�/�b��/���?�ַ"fd�Oi�Ź?<��>i�ەB�������	p�Qd����:u_��Q%�
%�~���վ���f�y1�s�b�cvS���z��:z�&���W��`���C�u1��݅%g�k��@�z���C7^�����*9Ti>�*=fѧO{��h
f��N]<oդ,߄��z[vPB�/l�ݔT9r^�.2%����	�N=_���Zhޞ[yF�Q(�%���c���o6�=5.[�ǂ�r����l�U���E`L�/�!f�l�o�����;TKU�����z��I@f�.k�z�(���Ck��;K�34��" �VY���v��4ɝq��,}e#�y���&s���'
6xKC�;����?��1���<W�q�$��V�j��mF\�ȩ��>ǐow����ь��R�����*��cI�Q�xH�ż�o������X����$�w����ګAW����nP؀��[�Df��@3T�잯�ɿk�=6J;�2�R�wy�TC�Z���W?��m��]��l#V�D&�j���A?�>���=mך���$�A�hА�� rp�D}�n)�<����łH�3PM�<ʔ݆�0S,��o� 8:�(\D�uS;/�[���k��{���A���s���,�v0]Ȣ}�bw��L��&���t�A�tSܷ�1h9�Hr�082�b	����k(_���YBZ�����1������'���p(ևm%�L^��.'RLS4��	�Q�i��@r#xY7��{܅.�II>��@�x*�#ρő��ĕ���n�'��8����/�as#�d'	�*x[���?wQ��X�Ɲ�#2l,X6���������Fi��������׌��[X�}T)�u��Gc��}�����Rw�s]T>wc/����j6�{.��k}�;�>/޷��Sd��'�{�t���O��ܵ0	�5���P'dku��ۜ*��Kkᥤ�Hg���9�� �����vڑ��MD�¬���/z�C̼9hbJV�XO4=SW�ϵ�V�(6�ۡ��-4��������Yr�����-�Q\Y���ƋUӂ ��z���՜�擙���t�չҮ��즃�����
���!F@&5-��9;)��\��x�[e# 3���X���#6v9h3��'�B�C��RK��tmG,��D0�dVK�ٸm��e\�ѝX�Up��ܯ5�Y�S�`��d^,�v���H�<�Z-���;�G�.?c����n��h̳�b1M�f�|�NoAv���0�`�W��V�����Vt��V��W;x2�=�vi��^�7_�Zn��ޏ�f�eg�o)��!�8'ڼ�0�X�|�A���~Z�h��I����{\��Ã'r�aE�T��%�R��LY�KY�TM��J��=����z�[�ui`��5������Qv��j=�	��Iʿ.�>������v��$� V3�u��� %}�N�D����X_���X�|�o�i:[f/��Q�O�܀�]@g	��tF�,��� �
qC\f�Ŭ<�[:>Nٲ[t�$��/����{VV�%+��%���Z^�oU��oB�^��)��b�M�UU,�����+��]�'5�%1rf���x�ĔR��[R%�F(Ƣ�� ZAU%�Q�~��2hn~{W�r/��7'�֫�������J:}���|���) Ό��9n2lT�y���[�:l�3�������-�4JE��P=+'�����l>��&��p��W'�lOM$q	+�X'���SZ���ug�΍	���ɐ4� E�X�dm<j3�z��)��_��>�?M>3�]+�z���b����%��R\�7͠n����~�0��*���`U���0�%ѝ:�U��K=i��~���y:Q�j�&=��qO����
�g��2�m0,�z/$I�Ա�G��GRآ���-Q�F�=[>��YFy��FCd@�-#����;~ �b���ч8�<e���X�q�P����nf�z��w޶��o���X���m��r�v�E��'���'ꆯZ1X�OM���>��/�Ȕ# �?g�����%�$4����q�oJ�3�ш$���z+Nz$+t��x�����l����ꕺ���w�Z�D�P����OR+�Z�GG����\X��f<aU��tQ�C�"��w:�$߷ /Q3@��D\H�s#��7����A�@����U���Pgm����r�@��+pbe���u���[��lYO�8"h��vj��}5"� �CnWC�.���J���%y�=�9>b�B�ѐɡ�+��g�B��x������ �,1�V�e�����#DPI=9����C�c#�Ӏ����	��=-3�N��L��~�G9n��P��,�T�3��k6�h zF��aW|�=�n�YW�Y��8�����9r-���y#�*͆��%X�.��0�ԓCF��<���x��t/L^��$o"-%(�!&�;��W�~�@��)� �0��y�0���·r��?�K��l?H�d\��x�٨��G#ۓ.��]S&��Ɍ�u���\�9�ܰ�]b]����Z7�X� �(o�m�:� �v�c"��]7��ِ�xu��:��2�Ε�5�ie��P�
-54 C�-�ŏɵRE,�F�`c���C�/�.�B.�!�5�Ċ���'��gv�
�v�u��+���
��W*-~Uf`��xϠ������qY
�����y ���j��
��h��X�G�������-Z<� �mX(I��NO]'P��C�~�+i*�q�:5�
�W��چwd�,�)�S��d��B ��f�����8�/�꫒HG�<�b}e�5�=&��~4��Q��},AՋ�[����m~4�)��0���
0KcQ�L����+�cH�s�X�r^߄f�#� \�3/�/����#k��	\��ɟ��,-{*��xQ>����!��1�� 6E�,a���ۜN�ũ����,�޽�{B�l�����<�ߖ��Ք�q��Jl��1���T:�L�?J��SG��$N"L�����>��^�������]�a�dִ,���tW���-���~!9(�r�~�t/X�MOu��((xi�p1����V &���x����q��k���%��MoHj�o���`a�3�����Df�;�/�q(J�:�򌍲�?9���"8���ac���?Cq�+����
��9"$���:>�Du�l���L��&���������	�8?�2���R�yL�GWB���P��~����)���B�	���	���t������
>�:�Ӯ�f���R�\c�����!�J]�˾8�@^L)��h��� 2��i���E?���M̕�/K�j�4w��Y
B�q(;kIb@J���e�3�����#a
|��FC��.���61�
�w�����eC~؊8��L���*g�L�>��4��ͩLq��ݝ��`��_5V���9���e��-�cM>�y�T?�T�^/���[f��jݿ�}�P�IY6� ��%XАX�km{�f��'��+��� �I|��L������]�}�l;��7L�_����q����?���E�`����Yn�,���6���sD��g��6��g�c�%��Fgz�$l��Y��l�q
���5G��˘TwX=oY���<Y��"^�.-�|;t����>������V��YV���|k҇P�r�F�C#�c���	��<����Z�
P,�ޏ2����Jk�������!I��,BB��A:��(ͼ������e�Y˗x;��ʂ����3�W t�&���>qh�,���[��$Dl���Ь[HÌ�J����*w����!׆�����7J&�@��I�����1{�th&6�X)m�Pc�k"�P�u����n^�q�?ؗ�6U�����Zv��ΥU��}��H3�����ȟ���61S[񟾷Mqw˪�����k�aVi 2P{(�[��U�̕z�.�� kV��s�:"��[w-C�,	�q�D�o��ܗ��͍	�4a�;�y��V��F�^���[D=�tl�j���t23r��M%𬻧:� >Jf�ۧ�x�!R���c�љ�'���8��_��?�z|cf�A���k���_�&к���_��n{.nC��Ռ{Z��P��zPT}J;9�p�</�a��J�R��ݐ�Ӧ7�#��)Y�q����&h=�iV�k�l�m3�c�Qq�pg*��y�t����^�^��.�/a�>iO���0y�	�5z�N6���@k��V��J�^n�_���(�֝F�t���w����sq����ȡ��~�T��Y.ϱa-Vԉ�Y w���;ѧ{>HI.�'<�U$���ɉ.Q��c?t��D�E֚ݯ�����ԍi�muz�X0�-a���յf�`��3F�Y�hʅ*�j-��^h��	<c@G$�#�嶉��&%��[�7SMK�a�4���ME�Z�����%����Tp�w$�O��EL
���L�"�!�>��
�d�Td"����㺠tV���JB�������6#˯0���
���J�M
O� �5���������i������}ʐ�БF/	v��uz��k
_�(�C��Q��(@����-���f�P�+F.W�����:��.,��,���YPK~�&��P�LjL����B%b푖?1�r��q��^�9�Fcl�R�R%s|a=�t�T����eFS޴ߜT&i���k�D��Nz������G�62U'��	%�9�'7��
��؋Bt�x�u�2��*�)�m9nr0_� @|��C  �#!ǿ�3U
�U^#�Bz��rRI����j����r�,�҇�U��cO�T�f�M+�] ���i��/����DS�@�7�kVy4�Di-k�i�}�;V�(-I�r��P�{C����H�e��sw!�G���!}Eb?O�����h�'Ǣ�tI���J%C&�B���� 1Η� !��ڼ���e�v(*��ϭ�?�A%Z��$7=n�a �6�%�J6m��}1�ѦN< Y�3���>��5X��;&Z6@јSu����ery�*� �d�^rE�EL�wo̔���b� �/�6+�+�Ղ�꼭]�	!vs�b}��d8kmVv)�eW\g��l�2w�&���j���Nx<:+)��)�y��#M�M�u��Ƽ�b���
X~QK��g����_~�`�w�����ypO�L��QD�#��ȔY
M�[�Eh�lCLCA�L��?n�ω'��]]3�����M<�N�TP6mh�R�����81�������Y��7��w��1�S�#�֮��(�H�8>�����w>/ɹ����jeڔ��4�Z�0mL�i�~s�3���ב�6#�Q���l<(l ����P'�e$��y�:箨����|��@}�>����b�TrT��ׇ��{�6�	ҿL�5K��&1vtZ�ϴ)��wn�k�+XRU:�M��59�IT�ZK�_���v�B|�z4� ��c�����k�P�����ֱ=!�J&hj���,�GA��*U��s]����.`G��F�v�{ 3ԷN�!��;�h�i^���)8f���Ƣ�K.�%��$E�١B~p�ξd岁�?�
M�-8o�&���Xr����f(9�*�6 /a�2I���>��q�X}W1Յ�����]ڭ	�}#tl"�d���wᤏ9�H�%�#�Z��$�կ���me�3ú��s�)�6D�Vҥx�h&i�iKx�ghpŒ�7�~��
||��f>6 ���ǌj�n��r]��/���^}�q�8�������%tU���V���,<f�"#8�0.�-�MD�x���t
��"� #�̐y�؈%� %l\�ړ�Pa`�����6V�ދ�3vB�X�p.�nI�I&�̡}�r�-�6k�*�i�\hR��G�)EY�Zv]�7�\� �=��v��;d�,�CˑWٴ6g'�*�ر����Fɏ]��(�:�T`� +�����s<&��c�-�B��ҹ�ަ���^�=}���?��KZ�*�I��y�;���IZ����K{~���� E|�.�@B�q�I)1o�2?(x&hN���e�(+x\����d��w�Kٙ3n����o�h���g�nX��*#��|%t��¢��&�Ǥ�h}��­5�gMu�1;e��:�(�F����"�ci���&P,0�5��s���ލӗ�h,��ң>�9Lשa`m��J7��0�d�h:��݁������Ñ����1��$���ONs�<���F�j��Sv����}��@V�;��i�F!ܒ��̬c���Xay�cN��� V��_,ջ���!O3��:R���%�a��<����?^Hh���pE���|Ö�g��(u ��q���]v"9�l�r�pX|sy�͝2Ot���g�F��h�ξ��|���AT ���D�1�D
q8")��/�����ա���M��9�&��2��k���4-Z�I��T����ǝ�Y���wōO��U?�ArQfh�ؽ���+hJ��:DV�}%fL���Id��^������J����
 �_��a֫��<S�$Ƶ���[:�N����׽��GX���=Je�7��ض�f���薠قmȲ"�b��ǽd�E-�UKoYA� �S�J����I5?��I$&F9A����5m5_\�d����[½N���fJ�3Be�7O[#��8�y 5Z$i�O0�2
�)K���i/8������}�PL=٢P�Tj���RnۋdjF����C�^��Z@ץ�[��A�e�/���A�)~�o:���>[���P�������F��<�J��q�fD	����'4�� ��^n�o��\����9��%N[z�C�$���e�x��5��5�6m*\��c�c��-�0m��g�+���A6��3���:��i�������ϥ���w�-˽��C�i8�SzK��n�/�n��)���-Tp��}n���(�5����G˶ ��!O�rwG�J@!���#�����4:�$A"xL��Pg��G�J�;۞�ؐB�<q]x��FE� .ߢ�C
)?J���%#��:>�ۆn� a���D3�B���nLz�^�L�JgՎ�v�ԃ�r�tW�Z�1����	��l}�ա�=5����0J]��8����r|6^��b��T2g� /خ�=�S��4no�	�V}��=M$!�d�J��.����<�B�*aY!Y�8[1�R,�@�U�fH���B��:��&@T�Oh\���Ze(��?<�{և=��-[���2�>��gk���{Ym�(�X@�B;ت����E}��1���P\&�\+������yT;S.tP_��fE�c�}y�B�L��m�nYi_��?E��mqEl:��*����Q�7l;���(jР�=b:���^7X�Lp%؉�wj�&���F]��+bH�ߪW�|��4rc�,S/=����M|�bf�UtQE�:t�au�L�AY�֞d����[G�^ΨX����w�a넼���W���c  �����2�nB��V�[���5���	��m�躢��L �ø�u��>��U�Q����ء�@�I~g�c,̞b�'[�	�n~�p�Caq���з�=��;ω�l������(�� "�N3��d-�����X�=A��$E�7w����2�I~B͋�5~w�C�"��*�j�ď�A
�>t\6-�^\�w��[���ŧ�O�iC�Q>G��f�N�n�vǔ,4��������c�(+�����&��0l��#���=�Z�x7?6}̉��8��DCDc�/s��*5_����h�qe�
�޿ܒ��G�������z��_0s��㮻�/f��U�a����۷ݎ�~d���"6~>y!�����2C �a��b2�K��1�WY�h��R���q�K�/���"e�Ь��t���19�+�<V$�읽��l05m���Ju[F��.���{F��V����Ѥ�*F۪��	�&�'T���e^,P�"�@��D��a,`\�0���w^����4��N�	���L�O��t;A�/�3�-��t� �^�c(�f�.�LJ<��m#�uQC��Q^ ��e��}1��S��n>��b�~⁝�A�7]ͻ�í��u��o�va�\kε�O3�:��x�K��|��>9�ÕY`+u��2�M�������黚��|&���5� �5�H��{��:Uf>U~�=bS�r��0�[=��LAz�J�N���~�Уfq?]�*ô���������z��}#�W�1@�M~���8�݅q�Ǯ�p��g�)C�<�]��l�!�|�p�f�?aĢ���e��tgk{��:)�QݻO�[�0
ǖ�a�
Չ�)qA��yn�/���r)o��?#��V*ǤG�M.x�4~��:a<�=�w�]/5"�}�#�=�R���$f���2��aŖqR�@+y<*�Ӕ��M-^6 ӈ�A���Iji�smƑ��T�<�n��J�Uf�~�3O:2HR�7#�����皩dLo�0�w��{�.¯.$O,6����ĭW�B�W:���|���[�?I@J)^e��f����������w<��P�Yk;�U#v7MB
P��z������t����T������npa�K|����s�o�<9��+[����y�}Q�g�:JI��lF	uy�X�2����"�?��\tS���b�IR�16G�7!�KeT	�'QH'�l� @��[�j��M?z-�N�8��'�L����̺�@�2d�p�}@��ҍP��5��];�����<-zW�D��:͝�e�a�g뼜�n��6h��iҡ��E�o�L\Q�#[m�51b��D=V�=��{Ҩ�@�t��M�������5$�죺z�����ٿ�/̞�@n�s>��ǐ)h �8PDw�Έ8��'M_ψ`�MS��V]�weغ��fF!V��\(d`P��"t�l�a�z�I�KM��UQ$@R/t'"V/��C ��h���Ex{377+k����9I���ȓ���pc���ff��෰�+�`l��$Kr���D�#�ׯ��=.ʩ���A��y�����Gp��7�O�;&y�2�2B<�!k7{���FؖH�˛-v繋K��}-�Үs�%�4��<lbь�vB/z�ѣʣh�=�lQ���=���U��H��EϚ��F�����j[pȳ��L!��2�V��7(O�q�%�Z?3��+.�P1��4d|ct���~f�	K(� )��'����M��sp���G���ިHZvєo郯Y�YOƹ\�s�IU�c"%W]tM"S̈3D]��)Gy��nF��c-�rRwX�h��%��9fAG��C��>0��ޭ�]>V�%��%��f�x�б�	��̧��}1H����r�f,0�����ì4q*�N+�0����p�S�f-qko������k�+����iZ:L@ u���_��K{�v�>_�/e�>z���)	����t��#�Jpӟ���0�o��ݍ���E��#k�&�}ZZ����h.$s%v�������˜�pK�V5;]e�Ȫ��P�{���i�tQ��.�ov�o^�X7��$�l�p�J�-�F�Z��r���O�dê9J�%�V��
YVc+��}���ލK�� ha9�+>���'�_�ٽo�^WlC��HAR�_�Fqz�
�����K$V�1W��]�%_����,.�f2e8*�@�4�R*�Ky��C>��qB8���� G�LiW�'^�[�}E�6���vg��K&M�[�C��͠�+�� >�H���x�\j�	cg/"��^�ظ 躺�V <Ώ��=���r0�P��=B'Ɔ�ΰ~%�+�l���5��љ3�"#��8p�1���h�GYpd?�=�\ju1#TYx{������zH2���5�+���@L�v���S@cݏqD�g��.w���Ȳ���W����:��D2�뤟!=�8�Ȟ�G=���-�U��4�d1)���J,�Y��w��$���BP�@J5�uJ�+ފe�����":�l*�rH���dv����"�l���%�'.2P��:��_�t�t%���R���a.��%}����lTS[]"�- �H���N�d`Wh��|�d]�4k71��ư�%�H���ς�<��o��Z�y˾�C6�e�A�${�֑����)k�"+��1��I�_�2#�����0���Vz�]��ᕱ���<��az�j��C<��渕�W�i�Jj�)�^�y�M�6�dy�zߦU��h���5}�9C:�8���6V��X����>�/� �虆�g!��j�&�ۃ��1���JjHvW��u6�9<� C�\lg!�`��&�����r:v4<���t/�^�����w�79�!���_��lq�A�vG�#��٬�"�"ϒ}H.�N�"�O��4�e�o�`�g�DF5Z_|����
�G��6�.��c����uz��[�3qv��(���`_�_�"�m߳&�V�]f���PF� Z�Ԭ��1��ܴ�ѲOɞ��ye{�eӰ*��0�헒����r�Q#9�&����Ia�����<��������SNb^���tM=cC/��a�ۤZ�a��ٌ�K���:���S�o[�Ӂ�Zv�w�-
ON2fH�l�"=���(�U[Nl֢k��s���W�1�-�-���D���#��Քg�Mg*B�D����:�(�r�*Pi� ��d�=���a���ln�ta��`^]�2ѩ�:eZJK U
��͉Mf];��[�v@=��M�;Y��#�k%��2j΂�b#�܏ET����U��A���in,�r��K�uȰz���.l;�L#���k7�{OKu+)�����j��F�sfCb �'N�_���k�0y'`�7�	�:�a��~gD�c=���81�`�f�n�Q?���!��@�`:�u(�6b��  �L�R�����|�A�Aq�/7&�;�(��D�}��|/�(�ԍQ�žP��K�EJJ��vۡa�F�ԥb�'g	�x7z	���$��<��J�]_��d�]�Q�E����d�w�4h����Qq.;�ys�d��]�.���?��t��;��T���a��Oj��~g�m�̯�a�b�U��d}��]?�y)�b��x� ������<%w��4��*�&��3�2Cԧ� 5�sZ�_�&�RV@���X�C�B����ˁ�2{��n��Rk���5��5���LO?_k4����u�y�͌�D�+������B�^���6P@0)�5&1��!������F%n���EN�=�g�d,L�>;s�J�m@`h\ޗG~�9Bf��(�ti��i��.��f��~��߽�+���i+��kZQǣj����u�`.���~�e}���MQv�r�V��G�oaH��r�f�"��V����!��n�+���n~TGM5c�}�oWx��2$1e m���ڤI�@Ms��f`28�t��i]|]\�2<�]$���d���͊�_�!���7y�o���e�Y��BkU���24%Ρ�K�"�ZE�V3������0b���_��$���~ePLj<�#��6(V/�ns$y'����q�j�5M�������E֖[�1���qk���$)��ٽAh���+WQ������&�MA�e"�Cʉ�d��R�e�X�	�m�t�X�m8�x�罫�ב\��?�3ڍ)f{*f�6�ԩ��%odI�y��dl}	���۔+1��)V����}\����p����%�+�?1� ���{I�R�H�*=��"&SZ�>�R���bK���Q_���{⋡�z�e��/��P�N��8$ �(�e�,J����y� �r��y��VPi�4 ����?�<z�)#`������(��c��U����L���G��k�nL̄+�r����s���H���L2��:R�2a�:O����'���њ�N]Q	�?@w�%��M��Z�uH�1Y��U�X�ے�hgӬ[[B��\eGEo�6L�~���s��Zrc���-��60�x�{a9 �L���h�q���?�gP�{��U�%AQ���F� #t�D(YYw����b�@#8�VA3/�,���>}�=w����sr��F��N!2�I*�1��U��j���K��&'2\����Ɉ��|���H����m6�U�=~����$M�j\tC:TZ����2�^�L���Mh>#�����F���2D�zh���.�a�'��ܖ�:4&���}ȔpfV��u� �!M����"�" �M�f�z����V?�kf3�DD�Y��t�$�F��Ԃ�?G�ߑ��=�.)�M����b�	�1 ft�2.�vM�P?
d�T����`���1���no�w�&�d���lvQo(�
��V� ����5L�.�t��)�;�V�v_�0(��*L7Ie��ۄ>�D���q��Б�����G��R�0�Βc6>eXb�Z��T较tp�y�� ����-�	^�!L�0���-����ay�B4��TO~>F����9.��IT�p��@	�t���x�;c�"$'y�ړOb%InTϐ���<�@���0�8�H���߁��!heD�]��k�V�V�"p���}6�h۾E���d�����J� �pc>?�/k�k��T�/�D�H�nH�YħK�K�9tt��.s�g�e��D�l���\����L�Gc��4OҚw�l�J�*0���  X?-J@N��� �]c��N����\ڞ�~e�	��=.\�
��*D=���eV�ӥ:�� 4��m�x�6��t̹���\)o��Z,�S�5��HN��k�_��~DEmg�#܀�aE�m�3�0薖����)x��=$������^۷z� ��蚉g)S���N��L+I��� ><·[�GL�
����TN�{W�be��������G�圎��'|���U"3K���SϽN@��Fy�t�;����\�SϏ���E}"����Bd����Ma6�/<��F�����~��!�����%���.\�0�Ƹ@(�r���	ߑ�+�6JM ��	~
�$Ǐ ���tҙ�6�G;]�=`W�C;ΦF]pR$�_��>��2�Q@��32�?����F�u�k���nZYH���k�������2�9A�����n>����Ke����Z�i\ ���J�5�Z~`^l��B[?�@pi�%f���C�/�W�_��6
�6�軲�j_u�P��Œx�f�9�D���V1��\�U�L��P� A�>��^r۹�t�Qhi(	[]N��v��D� ��њ(j� ��-?q�ql���9kS�
���e0�tf��h��Bb�C!��ia_v&�eS�/h}��UAcv}#0/�
(J�Ĥ��AVRH�v^���{��1���LK{r�/��;�Y�)�I,V-*Y�S*�F�2OD��q��C��Z�B�U����	�۞�w������
����Ţ,V���^�$���s�_�Y`K�Β:B�� N4�+b��M{��y\'�i՚�z��Yk��� >��A�	��`���m�JC5�Y՟4����{�����1���%�:�����+a9I	b�K-��ms�p����є���k�Ȝ"C���v��=��r����ǝ�2䑒<�I�PF�\�7'e��chaXF4)��_��äz�/^�V �/R��m99�0[F����f�f�t�r�Q5H�����?�nk��fN���
�\pչ:e�o�c��B��2|��#�'�l���[H��{QZ����MTT}�� �l�K"߈k�U?&��f�3P���릎�i�a�G�8�-֣���?n��-Qe�?p�I���o���Q�0��l�W����#�an ������l�'����@M�h4�O�:	T^� jE��+TxS��!�� �1DŖh5^L�?��<�f;~�G�%�|��
1ERҙb�a+Hب~��N`���f��nf!�'7�����<�l�9c��ݍd���uA�P��v���C��&D!����ݿ
��+��d>��d\�h���ԁ{:��u�lX}TU�a+�����&	:XޚšZ
��-�6��֑���9�7��@��A�Q� 5������ZQ2�p@�� ��{[��m�A�)Z�q1���¹�z5t���+�zZ%�a%�9H��I
 �$��U�F�e<$D+1�X0�4_����I��
��¶�9*�,��#���L��G6�Q����c�e��nZS����m����m�t� �Z�x��<�.���f�Ё�y�.^M]�s�W�,F�� �~pn�l��;I0Q��3�7�/�@�Z��TO�`��]����� ݺ��SL��$�{d�SG|���{]W�k����CxGH�2�b#*�N�	$�L�D�;�%���]�^��D�ϳ�h��zq?���aH׾��<�$�}�7?co����]�!��E����\��;ZЋo��
K�_��~��8>ѝ�)���C1�	���1[�l���ƺ�l��h������?�������(�8HF�c�NTݽ#��W��T=ER��G�B���i�d�ٲz:;�� �ǦU��$�2�/{v�FH��"�N�
�1�ǧ[���4���5ʸS���QQ?�_Ş��1�YwQp��^1�j[� G��[����=�?�A� =�gf��q|��קj��,r�@S�fU��>�4r���k<���nu<)b��WJa��L�L����Ui��_��2�w�"�)�;S��r�|c�n��:k�4�*X�"��g��^��H}[�q5A�	sN��+�Uc�Q��|��m�6�̏��y�j�rܞ7^$Y/���c)L/xZ:�^��:��M�W򀰗�4��{,�� C��.��~*��3W;��P3�z,\w�2��W{���T�D�At�P|�lL;�2Q�� �(՝���௤��CӻI��$=���E7���Ccd�vqu�+���&��+U��UyslĔsg"E�~�8��4�_�Wv�_���=�(,����ȱv#_}��a1��M���m�P�+�K��ϫlA�0��(�����Hq���-��G����Z�f�X�@�A�w��w�������n�e�_l�	y�C�������.���h��bZCL7�ߐN��BKD�<VE�Jɛ09;��k4�����X"{���Kqp*��xV�1��������VU����qk�[|�M�">���U�n���I�Jt����]x,�N6K筘0�:���I|��$1O��ّ`n<�:g+I�)H!`�N��g�O�_ �}HѤU�A'Ȯ	%0�Ɖ�9��n�P/)�S���NӽRg�t��cj %|,��NA�Il*��� ��4���o��B���~�*M0��D�~Ier+Pѭ��E�[�*bf11���.΂��F`%\��u~������x�����r�b���zST�㱖�Rms�4`��CkRo�[W��-����8,��';��P�gΠ ��1^�;�R�@1���7^|�z��!+Wo>��8r[9�=�a 9�tg�r)ա���A� ��*��Pv���)sʱK�B����?+���5YN�\R"ҏ2g������?�c�@��� ��СE�g��
�WYW�P)��w�k��,{��{��VD>W��o7�Afg.�u����V��nX�emy���\�T$�P��aFg.��| �?@l3eIU�����^bM9"����s��}�
+hS�x��U`}��mR�v��tB*��}zB\��e�nNp˹+Ό��u�o�K:F�����|Lr��W��3���U�h^te+�$3��Ov�U?��D��(��n7K���;X�K�d.֧B-0���
hQ�!U�U�B�]o�מd�X���0R���V�7b��3�:&��#b� ���cq?�/��5�(�a�U�� ����ZQ��M�ːL��(绎ԽscX���� ϱst�%�.�>��GR����Rb=i�R���6i����']1T\�<�@DZ�'�׬����{�|�ϊ.�+�������٩�$SA���jBF�D�_�㦢˭,^�uBWFcfM�ɹ�>7r���w��ܴr�&U�Xf;���H�4�t러<��� ��{M�Ak���t�Я�^��u���=��r
�Mg�7�� �+�+Z�o#'4��bs����_�V��7b�STf-�D�.�@|0$�2
A�M=�+����"�+��n�+�f��^t���Ɔ�H�^���~�	��3��v^d��"aH��A@ض� fp��`�^����y�ے��A�NꗓI��-�����EN�Jͭg�>)<N���w�Z������k�<�&��h�Π>���Lԙ����9p���Bb,(� �n׿:jP�ڽ�%��
߆��,yZ���7�}�E�uN��s�����ɠT���}f3��:C�BD���_����oU����m�9&���]�aT������e�Də�~�#���U�%&�v���Y:o��5��o`g^��ű��5V��t:\�-������e*�V�KNf+�33�@�e�H1�^rjA��(�=��!�`i��;�]�><)D�g��>��k�\����ʆ�,���Qq�9����\a��tb��p3_R����lm �:�� � �6?�-pG!�+�����[S��T�ڄ*���1z����ZX����S��Vg����#Ԣ��/W��h��@�K�z��"������嘈;?&'q�Bo���@q1i��2�S� '�"{ED]�w�E�W�
+[�������f�58y��Π,�w��/ǿg^�z��il�ƹ$��$ /�_QK�
��@�c�a�(��"gD"��H���l�{����Bd$���U��G�0ш�wG_�E��|��_<$��j�G��:CS�����.J�~��v�vt��,�Nl�%�Z�@�$�[�_��|�ڏ ��=G�V�ƄS�����h��D���6���~�5V�c4>�#|��6���`Z�c�����*Z�;�~�F���r�u�b�&UA��߀�R����|3�j��G�����49{��_��0c�Ud0/Ӵf�	rA�GB����4��(Woˋ�a��eЀxb^`a~~rg�}>�?��2*�R�jQLlx�9}�^�ᅱB����>sF�����T�NaW��"@ Mmy�Q�^nǁ�,�R��6���+�{�i��o��L� �����س^t�@�?*��	�x�\�jy��߷��ԣ̉��Qm:x�,`����J����C��ق���Ƞ���}+��ϭc����N����+"��H��liD!|���DJ�W��J;�r�&��Zq��j���fz��×�ϰ&��\_�A�H~Ri[R��xV�S`m���{�ԇ���X"s��0��K����+!���̜�
C}����z��@������r�C������zL����Ŵ+� Nda��n��W�� uV
u�}=�_�fht���.���"���n��~����+�R�	ި�@"��ù��ui���:�&6�ق�Aҋ@u0k�ρRY��ؼ6�dǗ�sw�Z
�G���T*
��G�E�6�ř�j�������tu9�����7ly#R�Oi�Wl`+8�����������}ľdq�43��e���C�~#eG:�&�EJ1-�c4I���Z5 _ʎ��ڍa�geSc@�P���-!p��,�"^d]�P:�Ҩqip�#rG+�=�_/qD�P/tCC���&|���m��䲻G4�l�p;���̇���rP����Y`���')�?��0�~�x+�R- �����T�[��P}���J����OPID�2`@��Tq��s1�a2\�I|���1�*�J�>~�5�ސi<5�fe"��P���ͳ#*��z�IIyw�QOr4�q�M�;��n�h�~��z��v�
H%��#O��7tK�x	7��H��-���N�i0�����M.h�X����nl�{N�-k��XEE~�m��JyW��.dC���_�w6�5�kBd�z�����r�~"��_&�3Z�*�'�^�}+��N��81I;�!Q���!�|E\�uc0|���1@]�H��÷����C�D�8+�_D�}��vx	Wk+(c�A)_�9%M*X����$��d ���[��3�p��i���K?ܧ�-<%��־�('�M�����|tË�#�����s��/\��ШV�1ZИo�C��q����TD�t9��?�����[�7󫝜�3t�������Ց�bV3Oj�@b��� ������:7���eЙ�/��%O�dcaĳ_9��c��%�`��Pc&S;Ɖ���T���7�o�=��cK:��b���ĕ�ΣX՟ 7u:kR�q�5E��Ҫ����`~+O�WnZ��{\��)�L�������|c\, `��޷CYCvɻ������ؔǕ��VS��F���`l�8)�G;���_5��t�h}��(�,Կ��o�b��Q�� �Pn�w�y9�!(���n�߲��H����#���
���y2��l����3VctM���1��n�p)������w�B�Υ�ܝU?�p�_�쟲��8v�� �e�ko��V��vh�B6L-���R6���� �q��.[g2���	oZe�'k��nN�gaJ����k�[{Ϻ\[�����R����ǈd�n�n��Y㷲�W���CKXC��*��0��P��#���<zgA�"	�w$E3y�T4��`vl붹A�G��p�T^ֱ���Y`
�����^r�
'K 3B��}�6 �z~��j.�v6��-G�]���&��86vdn��U�n�������䢙�����a{��U�U⠴Q$�v�-�.=���&�����_ ��־��%aġ�pt���!X�V13�aJ�<�X��=H���]:��`�?��k��BA��G���qc�c�VnkyAOl��R��ɏ����`�	ʲ\lp�f1,-�V\�܉t 'G߿t�!�u�V[ܤ*�7~�fOy0�������&J�����}��0�ab>-�C�ʂ�y
�xq�!�W'Q�;�v�y?�zv���U���y<��M(�539�ج��5d;�ޑ�"�T{j�7����t<�z�J?̊�ǹ��&�7��k���	e�C�c�E�����a�f6�iȰ��}��u{��M0���~�^#�� H�VAd>�[�5=[.��ƂP���2.STNzhq�����K�Ǹ��hXl�T�ObIp.��Lr#q(�+4�BH2�ёe<3���Р����oΐ�@<`���Hs�L�e㕇�zxK-^�MZ�`�ئ�:���x���//�b5�н-�\d�u���P��J���ж�%-�q�k��R)�ʹ!��,s���q��������q0Bȧ����{�d74�}ӥ�_��=����;����OX<KtYr	������Jl�F�NH� �+��S�_�G��H-�Sp'o��%?�wn[�='�%�I����K�m�-7h�p7Za�h#-���br,���5�%������rP;bE�i�Z�i����sg����Mi���`wN���3:�Ó�E�ʯ�EWT;\���d��v�}�~�c
d��).I#����7���f��D�yT\�1y���Z,����%@!V�����S�)	��qJ�>��T�55��'jEO1ԁY��a�_0~�/��%>h�����Y�4=�����d�Kg�\��z�+�/ʺ�&�kPޥ�4=G�'��|��[af����>B��8�:wU�{������ز��fV�!>�_©)%{|uf�����O�3 ���$E��v�_}�E�l^o�[�i�&���E	@�o�6�<*&���8��A�����`�U�gy�
V��#��q����k��h����&�g��C����ᰉ�痠�����4כT��Z�ʞ�8W\ !O]�/%R&�T>tұ����ǨS�ƽ�gd��lR��+����;H=h�����a��,�#�h���3�-�d���E�-e>}�D�mV_[��ʰ|��i�N�RV"��=���M���`�G&�(C.�j�<��k�"��S�>�����NUB��&�N��M���[WX�$6W�F�����T3/���"Ǐi�1� �-45���Y��V�[+�.��S0.���8��u+V���G���jv���G�\$���"�Np:�/�� lxT���P�_y�F�[�M����MapJ��_O��C�{/|��r��XA(���1|�y͹诺a:�F� =W�|f�!��X�)sa�2�>��-��O�׳I�0S���fb`xi+��}���0p��B������}�FO�X?��p�"@]H^5�%��V�-��r�2�#A��� ��,���k���gr�>J�������qٔ��2�5�p�rz��k����q��{��e��r��f0���7��?Q��J�z�؃� �E><��j"����P*�C��'���ǚ�JGL�g�4]|�����/%��
p4/�>+�s9�і�Xh��>��EZ�I��y
2��u�)\=���(��{Ǘ�3bПٯIZ ~C�wP�fV9���U�|�/[�!}�u�9���xf/�r��FF��
CWm<=�u7�����q�(���0�/��\g�F��.��ֹ��3I�dL�����u���g�5'����y��f-�cII��D

�(jh�����sY[V�`pS��ו�m"�ج�;���I���Ч������Q�9�y��6����"�
�1k;���иE�l\���M���$+w)��LAW����������k;f�+�M�p�_��01�:;:�z`�&�Ɯh�3�q�w���ʯLg��D�uzo������o�7Zh�����+T��Ɍ�u��+I�����O�3'��KCpIY3�aF���td�ģ@ϖ!Z�4c5V�"DZ;���c�W����I6�^P��O@�&��q#Lf�\b�����c#ǟ�7�Ơ��縞|�9]���}7�;JH=TB���(���-��z�G_f�4Ǆ'#�T��� ,��Ý� _ �㘝*9�>8����j?���*GN���O#ˉe-��V^�I�t7:��C�����Lh�D�U�\[�\�B�I��~ł6�����C��4�#G9�9���r�6DQ��H�;����L@�W��\��<�X���}K���X��a�A��w�A�	���^0Ɵ0��pZ���*������9�_��>ݧp��@�zs?d:�?xP������Lf��tW���K`N�%��#ѣo4���Ō���� ���{��J�Y�ۗ@��'������ڛ��[$'*q|H-�]^K����rı�٘�J�i���Wqˑz�b�LEJ.�Χ!������� Q6��p�3\�����1֪��� �����lq�J�g�?B=�֭нVE��O�?m�c�E^�	�Z<��Hߍ��o%��Ĉ3�u�-�a�H����h �@�Dƈ21Fm�m_�Cp��ڮ�B�����Sjd+��$^�=��d]Ѭ��7�b��)�=���α�\4}V�He �4�a���x5Є��H
!���TM,�o���:����&�֗�v�'k���=6=������^�������g��1G
P���ڳ��&�{�J����"�$�3�>�]M��y�x.�,؊��˓H��JMFi]��74/M�-<��d�^�o�-���v%WM����x��f��[GD	���ޛRK������a��/����=��o��.b?@Ҏ��J�j����e��}����K!��̃�� ���F���C�R�S'����px(��;,���)E
`,��h�/��z�A^ �����8�����v�[hzxc�C�zw�U�gL�&��c���$nS���{�U�IO[��"J��F� ���!+i�ԽC5��4>۟���?K�\��YnK�*�7�F��*:�
�� ��L��k�K~M_�J��������wj_��PXŜ$��yZ͇�e�c�N�p�D�uD�%�!�	��W%����î���~@�����;C��~�`�A�Q|��P6���Pإ'G��G�2�x3��p�����yV�$�F�C��^�,p>��7�H���8��ެ�h�c�_�g�+hXz�z�C�y��@,G�3?��X�8�#〘�F�4t����W �jK��z�!N1= ���`}ڊg�}�Q��F��Ofxq.�|�$��ჵ���ŃN��0���?�#�ߴ�bmܨtz!�VK;�9��GhcN��z�y�!1��m?(=��g`�9<KC(�Ɏ[��v��`Qr>�>R�!s���DY���E[����~-�8�!-\�kɸ��O7v�bt�S?�ⱏ.��_%YOȫ�S�`eO�埒ٷb J��6�$�r��K� 씯���2@X!I5�6��O�M{�+Z�q�a��l�(Fx*z�,GE�@��8QǄx(e\�B%�,����G��ዓ�P�_k:�4���h�$cۉe?�	b��V-�=��㭨!��\���S�������U,,uX����H�����>^g&�w���b��;�<km�ϩ6å4K����ýTۊH0R����H��rk4�' �\�w� �	t{��.�JF�x���kƕ�%��-K��jXi��M����D��̲�d�. A,����<��=(iu'�M����>��j��I��h 3��E�ٸ�=vN ���'z�C��֘��z���Ne4��D�����Э�7��������[�6�olws2u���6���O�2�K�H8@=�KmK�|[�0�F2y�8����$J�c�Ф��P�_s�+3��"��u�A� ��A�5"o��wn��I�*1aT�t�3Y��/���C�����2�$����x̠��~�V;2m�գFz[7������ga
W��}��n���@����xe8�V��0	릗S�R�N�Y�U������tl����@�Ώ��$K��4LT�ó+b�3O����` �׸^=üi�B �]Sss�HY�i�x��#���n�E�!+�;?$�V[[�I.L����V�H<�QK�1��`�q��*��\"�?>���=�Y-�R�e$l�4;"r�7e�'��}H� ��T=A����;���G�����}��)��r^�-j(���wqS���GrKc�ٻ�`~֜�qm�W{��ёz,H>��ՠw�ޛ� ����7�5Y�>�p4ԅj��ߪ��T���u�_M^<��{��r��`���D[9{\��:�?7.q�P�g�:�<k��}��gڹ�Z\W��P����:������b�D��~��Y�E��c����M�y6���ǻ�ь�Gw82�s�J�C:{hR��jc���&^�` ׽3��Hf�$8y5�J?��vYD%�D{�/h���h��ItN�=�#w{�*�.,�X��W�U�6@��w�h��_}fP��޶;���eI �Rt�SP�&��@�{�I㻣�>�\��#�F��OUv�J<Ӽ�����B~ll��is{��XW�D����_��B�@�1~֘������9�~�������|�͖:�i���e�I��ک����3��	0X:S��
������{82|7ĳ#�����(�}j�T�<p6$?��������j+�_����C����뽡2�ݟ�V������`(M@tM&�DL��~�����xo�M�l򕹊��Ɂ�Bp�Xm�O��!"5��ZՂVP�(��:CQc�9���(����k̴{�,t*"�L� 풱�}b؛\�\����*Q �y���L���'�%�k�K$�~���p���q���:����-�fn_\���P�S��m�1�vl�&$iL�Ԫ���q��4v��/��Z���*z�  9����'w�Ȏ�)�~
����!�â���M�5��$ЃA�jg��"Ʋ����d�2k؆[+1��O�ZYT.�ͷ%�OXC+2
�o��5�w��X���� Xy��cr2m�p�o <z��^f�ɧ3
n1;'�`�i����"bԦ�l�ҏ�U.��E�J� �h\H�֒�������l�� *��V�dvT�?u1��%�]ٛ�21���.�2J�6��s�s���zO��J܏���zbav�m�~3^��W��eUɽG�<	E�m��������
�58���#�r�b��ց�A?��^�w��;/��zF���|��V�:	�L=��k��߮�"�(Z�5�\���M�� ����,�P�woxx�逄�5�A��~JEH������^x���Υ�	�cD@.��ps�¦hB���n�F��I�r��aͣ�m�$�ݤp|�Ϭz��1=T<���Fop�C���D������w@u,?�b���ķ�>_�=��v�d�F��
HH�{��	�3J��,뮮��?��C܎}�mi�7��eor�BB�$楯`��Q���'bh��K�=4�Y��i �� �����>ο[�ofz���|z ���#E�?�ʪ��{�N��K�c3X��T�:�i6E���FI�RY��5�����UY��1��EM@��x d���K5f@J�N��.�Dn�t~����!��������V�n�U�`
}���%��!�M�f��@AK�Ӗ��@�ѧb��(B۸O�j1�['.���l�]�s�;H_�E�A"�-2w����~\GP/�d,�/B�����@��\q!�=�<ѷXJey;�a}<-a_����Ȑ8��;�#����Q�g�q��=�'8n}]�������B�-��b��?��k6��Q{d�ݔu����pF���U<����3���#��i���S����\aGR{`~���#V�H���Ty�*'ƅ<�B��i�X��Y���V3�`KfrS9��&��
v��U2���/��'f��JR����z�A�s)�%�+��Z���3�*�0�q\�BNx��V1��@x�/��k�k��$��u���p�[��O��(�鑂�!��c�駖�Ix���$�Hhc��$��?���J�?��D�ߝ��"��G��jD$W�$�ю�h�uu�`�z�Eޔ t��+��~T=m!������YH�+M��|�Ϛ�3�'|tOTE��KT����xnM��h�NXs��['��D3�d�L���HZ[��A��V^�3�C���a�鮝�<*QN�s�������O?w�Pb�{5a�����u��ƁSM�z��v�B�	�]�bD�8b��m{�9��!枿��873͖��z�Y!j��Y�^;f�>~]�.�R���,���_��9�U*�a�ʤ��Rp��M��s��g*ѷ�MS3�u&߶�j�[�S��dI��j�<���Ϯ̘6���5�Dp_�ck{"�<"��K7��{D���hm� ��:� �#�Cz���>�����H+A?�V��]��$6�ύc>� �
M�.��ml:_@2���z�ݥ�v�$#����z���'�:F������¦����||�c@������VR�"�j�b�"������w�+䎾k+��rt�9�~\���k����0&� �<��?�7c?/�Nz4��/�w3��^w�ٸߌ�eX2��a6����j`��=�X�-����u#�Xh�`p��V[(����m>Dq#� �����TS��/�W�ЊΌ7+J��Y�}b�ڕu`��h�0yoA>��f�_ڴ�߹��߫>�m(m�l�4����y>���*���|����F��PSnQ�e��������
4|��\�?ܙ���N�Q;r�ZDԾ.C�y�P,��Z�[���(c�2 �H���^�e"h<x��m��2H�(U}��c�
�M�
(@��M&j9��x�7�@����uN�!�sBH�A��B�`F���¼�����<�y���+9�^0� �la9=�M��AS�1  �8�좳�x�K���z9������ �w�%�>3��J�B�3�0r����M��ZCE%տi�.T��(��,������*C���Le:��t?#�H��h��kc'q�	�'�
�M	o徒y�)�/����:T�9�c�ΛӒ<�{���pA-;��ڰ;�tZ?(:��Z��+U*�U�6qZ�QyH	N�]�MƔ�b�/n��#�(��{�0�����8�5�-�ZO�lQh�ƾ���L���;j:��鯤 ��Nl��:�4A6�x����~؄>,���7$���,c
E'�M{�R)��F������2�mxJf}:�-��E\��\t��Z��0L�g`G �]�De�`�{���i��j̆�z?|ʺt����:��y3��%�6~���]�m��=f��;�2�IOӵ��nb&��)P�T���<2N�I�*�;K���%ցR�o|���������-A?��m��ud�Q�N\%)$���$����7`^���"rR�+��gp��&=J_�^]`. g2{���7e�Q��#��h��O�W��m@�l�ff�{��L:�H^���8��$D�1@z���Tu8�T[��#
g(��[�
q��$Z��%�3 ԛ����b�����"�ܾ^ Y?��-��;Y�e��n!�^y��_�7h@�h��%�����:�.�ښ{��{ʘ^��D┰���8�p���(oD�g42</����7�\`���T�>Qh�������"��c.$ZQ�-�d�w$��wls3;���آ8t�;q����]���{<��R�m�QeQ�9�ӥ��Ό|�Ê	g��Oȱ\g��oz�QE�$��1���;��у�:�m����=�<|�� \��"8�����R��"3q=��U{��w;�']�y�� k��#'���4]��4_�\r�^2%�p����p� �!@�GE�w�sm�8�Ú~���Ճ�f��̍O��~j��z�o�����ވ����Ԟ�O��O�qU�"s��C7�KGľ�:��A&7��̔���N|�;9�I���D�w��W6߳ >�̶�f3i��ah�W/���H�`*���/;Z����/�Zk�����}��֮�Q6?�K��Q���hA��fk�VGƐq�N��Tb׸"������+7�"[�����%����|����O�*لf�G�3��z?:{�D�����?�7i�sK��Ȼ>����;JE�(Bu��l	q�d��O7U���1��f3����L��U|?%�V��}�i���	z!�H��V����QU=�>7嚾_�P���1�Q��d|,�6�]��zg�c�Sp�w��.n0uz�ɦ��qu�.�/�����	�[�(TOo����������h��@2L�)648I�M��YZ3�%E�����(b���]�7����%s�����#D�W�]��\�m~$�^Ygr�1�g���8h��T_O�N�i:LH��;���J!b2��x�'�&��\ țhqC��>N�����+���a��N(����Ӫ�ApU��X�t��Tb���,�|���{:T�e�y�2�1�{�5Z~�Q�̍�=|���4�m�˩�?9�@D�g��f���Z���m�m�T�<?�9�x�R�r�Z�U�r'C5�����1���!��wc�°a��M0>I�+�W��>�D��i�/W#�����ޫ��SC��@͇M��0�.�*�`db�U#�oU��ƶaA��@w�S�J��3��
}����m�1_E��T%�~��Cƭ6��;��tٛ||���n��#���\��jGL#��[:T�Ē`�ޱ�)�E�8]��4���(�v��,�3�����^���C�R��!va Ԥl�.�.�}��2��|rS��Õ�G	T���)F���d�f��`_�dE'���6V� s��EA��L2��I�[ʬ��wo��m,�8��U�}ep�o�ou��گt��S��Ӄa��ګa���ĸ��#�ڂ���
��Vtw��_[�����?q־�'T*�k�{0i����SpP_'9ܠ��_z�GJ�����3���|u�V�vvk �*�:�:5���9~�09��%h qt�	�����r�[��{5���p����|ܱ�'��*�Z�sH�XP�F񆷆��J!��#�BM��;u�� �fXɐ��᣼<�T9sM�Bt]�?eZ�{�^�jE�k��]��P�^�~}����= ��̝����&����׵_�z0�t�'iS<ctq�?���.r	¡��];a=>nĳ��#Ou*5A�Z9�(�\�&����.�n��`¸}Ы�ǘ �G���lNű[�9�(0lެĀ��Դt�����І4|�>�.^����(k��~o�f��:��oA`t3�ˉt�7Ķ�Q�a4.�*�'��3��X�f}�)���">�,�� 0���p�B��D�ϰn]�9�jf�<��}��H��TLc�(V ��Q���~)ؑW�XC�a潦�m͑�v"��Y<�����y�����9Ű�*�&�T��t	}&Qّ��}�P��ǂN�/��tq�$��+�z"�a�GЖ��`tUaʦ��KS΂�^Vl����թ;>�`Xþ�M�E�Q�(�=���pTf���V�!a|�d#]���fA���抶���~&ŹY��Ԑ�	CϷ�DZ..J�\�]֢��#ރ�J��qǏł�k(ȾF�Iܬ"���L��D��p���Ozw�WUԯ&I�ః|ގ�e�z7���{io�"2�l��K�y^
����(q~*WU��K��
q������'t�{�$g�C�Z���E������0�S������u>L>?�l����R���뢇g�T�IYo2�R�-'j&^aL�XwN���ܦd���לA��N�	Ѕ��iǪʸĺ/g��ȭ���jl�T8���v����񗽻��#D	L�"�(�=��JB�!7�z��r�))9ǘP�6~�|{O����]���P3g���v��)b}�v\�r�纸?�i�&c'�F��Ɏ�Ӡ�9pD"���[��ײ��s��i+ˍ1Y�r�U<%�U��Z]��Ügc�(���_��-�d��q	#�ɡ�ڱc��u���Η���Ӫ�zς����ZY���i����=�LI��?ǻX�5H^�b(�QT- N���!�ZƑv�&�\?˾��qɱ��R	F �ҽ��,!��p���r�0����?4H<���L
 "�_ �7�pJ�kr6X�2�|Ȥ���xk��9E-~?�0�<����%c��eq�h���u<&ũLӈ�Q�!���s�����G�`e_�!��6�;29��t"KHy��>d�E�Q���@�wP��|'�zM�~ڬxJ{�A�?�+��,�~�x�g�#
�7F��S�@*�3��$�`f�}O��n�X=bդ]O	���7��A�,S%TQ�e��oK���#&���fڌ�O��¹V9��4_6C��B�����&@[�ՇJ�A=�yw��|����9>��os�c��=����� �4�fn��Q�On��eT�AE(����H�.R��!%����$�`�鯍{�[����G��E�����b}6Vy�tS/���y�͍��Kۘ<����-ɐ���G
.Z��୴��ډ(�D����̼?�w�Bác]`W��R�r�	�@D��%!���<vh�ŵ��]"��|���J�����FS7�H��A�%%7�l�Ga�.���~M��D�\CJ��"'Ǫ|b�a��S̏
B�~ф�Y��h�y���΃�#���иH9맚���І3��>NĿ� �x��D���|�����)0P�7ڴa"������|
U�_��-�񀲩���L���u*�G�QRD�"�"���4��r�7٠�X��^���Gz����c{c�5��ɾ��R��,\��w� �Ӹ8ǈ��B�t_�MA=�Ah� x�\��|E!'��$t�qBrj�(K���f9N[�q����N{�-�G�Aׂʮ������d���&��ů��T~"�VJ��?�ρ�j��i�|�J����A�� �?;^;�k��/vz��Z�����#��I�m���D*�͖J��=��6-b��Ӥ�'�&����0�q�+l�Q^�A��}V�6�ݱU�mۧ��|����B�8}ɗ5d���(��8W�����$w�%*�%N�Ǡو�y>��@��i�v-�2�<�n���6���qs�����
P:�������T���RZ�P��2���Vk7�O<�5M��`4R=�#_	m*wK�%��X;%G��5|�j�	J��1K���:[�Y���ʂ9��Kͷ�yM<:p�W�rWb�l�Z�:��1�ఋ`�h�:)�/^5�,]�� ���Ò+D��EL��y���З�������ջ@q;M9Q�����������r�^�_o��y�4�N4�-�bK���`S��U�H����5*Gr�#�f�$=�	���?��H�ҹ��ՊT����*�����8s��l�o�Aj���@0<��W;��h��U��*��?ҕ�FU>�S�g�!�g��%��  Gz�	Hg��}��!�췰�,�7�OO/���V'y"�Ku5�o���k+W���l�+��_ �5��kV>�B��mxB
j qWI����h�#���EB�#���ē/i��9̖��>xt�?���(�PJ�,����F~]αS!�gW�"w �-�,�s�s��~���P����l6������?-�jH�0�ի�I�;o�u�k�7���2ѝ��iq�nTL�mj;L���S�V��4�����hBJ�"�=&g�CY3�JH�0�0�L1�}Mm�/�np�z�oҖ��f z{V�8Q|j�^��#ɒT�R=���k���v�A��	9%�Ez�Q!1f#��o�Ae=?w�������j[�c���H�(�J�a<����I��p&�����hw��I�V8�)���E�����+��o��r�&��Ж}������}*9z�0&u�G�\�"5Ig��,B�p�����$��[��J�D�
����(���-��߂�PJ��{�K�%�I�&��$�������tsDC�zG`Y�+��j�>G�V~ �#�#H? �!Ȑ룄Gr)���o���0�f>_��_��k��.l�&!�v&Z��C��E)���/�ZP��k1�b��{�G*-!�r��y�k�2H����B$�k���~g)C��8��Üar��%�)tggi�r���X�ǚ���2B�Y���o�W�un�-��R1,���a��P&���B�g��h��_c�o`]��9��Bڛ���T�IgW�U��z�@�7|�*��3��È�}����{6��{`���+���	@�!Ex�<~%ߪ!�/����^����`��`���}��0 ^�o�ǫv�����V5�L��ΗVCJ��Y�Ӆ(����a�,C.k�`�+h��ٝ�Ӳ`1���oz��$�GJ�Rb����v�*�W�������m��m]�7U�i�B�s�<?��20�,$sZ"�]�LWd�h����	��h����U�)x~��j#�� ����/�
�GX�w�wCsY�V��%.�kXI3I���YuU~|�{��<�yomA�o��1y<E{��y����ȹ/,���66E?�M1NlZ^j6@�� ������=�sCf�Λ����A�03���^%Gő�g)��n2I�d�ӎ��s3��.u\��4��O(�܂���9h����A�kS�1�*�7�5�7�m%U%�8�΋���'��L��;���G+3�2_�\������'�b�`06��ڜ�)�{?��
R:>Y2���*m��ZfD�r)� ӗ�FIj�fw��<�3�ⲙ��(��4ϡ�8���a�	gӷ!��	??.�L#
dj d�wѯP�7�E���Ր<ƏUw�ulg�4�D:��z��4ŚЗ��ύ�Ӕ��u{��Ɋ��}pZfˮ�r&C-�F��꒗&���j�uI!"Sq���bhC5��_�vg&SED�(�g��T��w0%��ݩ&XiK�VR����2��Uy���k�t���������M�̚w��~�~�|7���ۇ���C���cy����r�
��6�"�b���$�ڏ�L_W�Pf ��-(�T������P��%s~]����}.pD���Ή��d3@�K�ï����`p�3��(�gN�S|��_�RYSn N����i@�oΎ��N�è{��l���[]v�&��q��~^��d�ײ�l�v�����Z��g\�կ'�-d,Z�8��$��>h�r&c���X���U(�ٲv����������[�}�gMtj�BcF�l�x�ZX��^|�����T���D\-�˯`�\�c�8X�Нqh�5�D�6R�����%(��eh0��X�) w�����F�iXg=���0�@�ͼ\��[A��u[�p��J:�\�^7E��Y�p��P�s"�g~btEL��@�ee�7�feӼ<}��r��*/�gTeU��|r�X�]z��*��༦5/u�����l���*��#v�F2VV�2��%��m=f��]�^��%����/slu�H��E
x�%�����3Rhk%M�^�aK�A�82Q�7�MȅUڿǯG�I(ὸ�'B�k�U�F,iE��LI�cS�❽U�������n�9����y&����WJ+��T��A4��#i�8�PUUI��#��A$�M�}#�� ^Z�ؔ���뤳�E�Ǚ�P�����'�C�n�s��AzN6�A|P�bH���|&��K�Vw���)E�8�%�'�;��a�YZbU�kM_X�-�[Yv)|�>W�2�����%�j���v6S~���=.0�����;���zv��V�X=�M����W=Oވf	��������ĕ��-w5��s\�7nGj�stD�<�0-�K��$eWΈ�p-�îl�+�]��<�˯�R;<��yc�����lH׼�T-��c��Ϸ1=�{6_���K��>A�i���"l9@�L��V��ad~���Z�;;���\/����a����7��gЄv�a����� ���XZY"���_��$q��������N�Y/���KV&��mJ��2�'7}u�7�ϖ*RGR5SK�����^
D}�&!��h�咾pG���o�<<2�F�m
�qY�CZ�7�?��a� ���u��s���d#"�+@ ���+S��|_c*�bV���~VF4���	3������l�<!��,c@Zt�n0���BX�y���Sz�L�����K��Ua����n�s�n�D�ct���^�.�?r��7B��8-^y>i|QU��"%w�x���|9"��L��y���4�C$�q�?$8��'�p�>]��]R�ʎ�=��[!$P$��i��^(+gl���%���3IZ� t:�&������Y#'��"bȴ&E�Y�DON��tP#uS�%D��Ղ�Ǧ$ͭ����1���.J�'x3���?ʦ^1|��M���$'���G�KF(�Ι�n���˧n��A��;ܭ{��ԕ�gQm�+�t�:�UQH�fN���V���!>�s0�����C��Z}�1f��M�H�����4/��ln����8��I~�*�H?��ɘp��&2y�[ WNa�u�9ُ�K�C�p,�q��$ꀸ'aVۗB��$�6b½�q�Z�@��7�~Q�)!�k�����|�/�uA5;A)��u���veĉ).b��^e�xC̊�r�h�&AaBϚ�Bi����=
�p̺A���ߌN@n���H]��4X�Yʱ^'}�#�k�m'��Rǻ�-�4J\�F���aeA}�r�U5=|���Ϛ�Ƥ�j㬵������
��'�~��t������I&�>^��9I-p�t�y\5Q�'��|��/SiQq.�+��>'��� Y��c� h����^��2Z�Wu��!
<~��w��݅�Lyk�;U����耇�N�r,��f���x�-�̪��V�dZ
Y���EB���$���j��f��`{���Io^�?,����S}r��p��񫜊�gG�2r��tXC��_.�0���	ںKƮ��&���x������O5r��">��X���"=B��	��wU�>�bC5Yv��B��9�,��"L���0l��0$���;�u�?*ʿo~�� Gj�
3� &0��}Jh�2���}Q#G��#�����ur����vv�ǣ��vVqL��GFZSj���x$ZF`t7U�7G҅�{��ӵ5�u��EG�*&H~�h5Y����S��%4ʣvkꃸ0cWP97��٣�
!�E�PK�lyN�o)����\�p_\�/��&^��d�#0���	���*_����t��7	����!��]¶�����o�WH�o��J%(x��6ha����������"�sLڸ/R�6�|�a8����ҍ��1�س��~���[�&{�c����	yx�B�	��K�

ҷ��2���q��=O��Wdi�$#��.� ��}�*,�;���߉�"���1 8���{!�4�AP�F�ӽ��k����)Kp���f<����o�
�!C@ć�FLr�^�W����G_��A5y���iL� Wj���<�%��(���L�%��+��B�to!$}�{�)�M������y�rD67�t��f�w՜����1_w�l}�V�md��1�+�gi7���-������]Q	��?]���	ٳ�GЁd��\�-���p�����~k�"\g�8�yshӺ�����D��[&�3"���T�){��V���U9�q��1Sr��^�%@>W��2��c�M���Fe�dϪ
�g�jEt��Wb��{F�T�VSf�<���g������%H��H^	�Z��`/�w�
��}j=�`,�`�]�<@��e˻ۏ�X����o�ǭ���ߕJ�+��;1�pQ涄�˪����a$�tD2->Ĺ2�5'T�r�2��}�"x���7�cP{��ey5�L��$�S@��	�k	}`+�	���\�r���hך��_�̯�6]��}p^-�O_�?V¼�N�� ��=�Y��
 �ڂZ�ҚP�Z�>�k?05~�[���N��\-ȯ���.��� �GN¤(?GLkǦ0�����,��)6*��}��)����#hU<s��d��yBڊ0�teu|�Vz�4(ɒ�FuCށI��έ�GK��VE��j]/�$���>
Q�@B��(�2{��*V�V`rgjAXգ�y�P^|��YK\�t\��K���lv?�*�Ǫp]r���e�Ǝ�Vm�8�f�_�6?%����U�g�3��N���sU��-����:\n]��="��/+��|��9:O��Ud�q��١χ���[Q�ͺ(����`-1�	����2t�3��t�)��@����bj���7@Kb����צ�u���B���	���#8��'w� ���UZ�U��O�[�MH��3>G[P�^ܾv��|�Ҿ��ƪ�o�gX������gq������Kڇ]������ ��gx"L|D�����fxmJ)�-h/��O��OՒ�E�nȸ����'�.�rv��h��s��<X�˕$���h�:�xS�9�Dg�b[2(>1����u=�ܙ��� �z���M�:��L���2��� 1I�WҾ�K냵QD�E�l�0�4�qϜ���t=��~�m:d�X3I1zƻS���SV���^�@����4]/a�QS34;����Ԍٽ�&�H5��[BwP�e�&�Qh�_|�54�c�5kB��(}H�- 4L���ϰ��R�<�x��dKX`!p� �YFє��e��~3�.����T2f����_b�W��w���Ņ��֜��*��� �H�g��
� �x*W���I�h�VT�B�G(rB��z���8X�I�f���$ �H/�ߢ�h��j��!8�[ೡŞ�+����b]C��رŋሂ� ��&)5���[���;a2�9w*��ҍ��>�(���.��.d݌P�]�埗,W�Yk��CMu;E��s_�R��A�[Z���mM�|
�}�8�{�6`�dƅ�f<��E��"�1�֐A'*��g^v�0}�G�W`�������2���e���(��O�?��>����ުڸ&���N�0�t�r24�3j��l�{@j�p�L��k�v�C�b�`��nϿ��Tn�1�y�O�
�:���K�9#=�C��B��K�L���G$c�@">Ez�O�<��Ԙ�ʬe����}h��l
�(�ע_��_��i�Y�B:�y�Eɝ.	�J�D�c�����t�u��DoB�I)��	x���ΞH[EΣ. /f�v�V%C��2�y�JD��/�K�~�+yH�f#QM���ǜ^�.v�ԭ":�{���v:n��DȨ��L����9�&���}�P�����"sy��Ř޾�?E?�$������&���#��Yt^���l�m�Ӈ�2�[I���b{��AB�[2��\��/��(��2G�
�Y!�5HI?:�{��[^��v��it��4 {`$be�5u�)##6OX`}WU/L�j�CZ�/mm�c_���ػ��T"w9;�� w�?�^:QzY��	4�s����Q���C�b�k*��T�iEg�ް1��+�!v������Q(^��Vb$��!��O!��<n���N/��Ӯ����nTY.Լؒ�i?l��� �m"�	��/��n�����qd�{�U$1*'�:�������&��!?�qt�R6,&{�p7e�,0��k��}�%1B�8�>�Κ��u�X�,d{�+2̍@C�;��d.�kb/��8��4s�v(m��hOWgE~��ۜ򸆑�Y��N�A��,U9J��1��E�9	}�����F�����ݽ��l�{��'�D���8�	��l{�L|�^�o"�~�'Yl�:X���s�w���:l`���Pө��0R�m��J��=�����=��'#`�6�d��/�4�9I`�{aLp���ㄝc��MA�}m�2�q��H�v
�{�c�;}��=��o��'ڼ��	Pt�;����Vs��#r>�x\�5��f[H%$�=뻐@)lx8`X[�+�:���A��:S�����ךԎ��K�w�
��/l^��(Z�eg�ǄU��y�։�����K����
��T�uz��\v��wNc�c�z ��L����>�L�F˷7���ϋ2��3���Ng^H��JɆF	��}J���42��L�H�eB7�[�G�%,�����@����b�&8�l���Ǡ�Ű�!��v��W���5V5��ۇ�$�G+�os�.y���u��;��@`<p6�1�1?½R;y(I	��2oQ@<ƹr/˩�g�Q�����&=��g��E@�e�cY檻ԕ.f�Dߖ�&��?^�<?u|��==����]Iǃ�_{���#�������.�Xz�Vg�V$gӨ���x�����-�n<�ѝ��y�m��KA`�N&��v��O.�үpc�F{����4c۶���=\�����r��D�M�����y�e���MkE�7����4ٖ�p����C=#��=lc�;?��_�wh�_P?��6�w@���|aK���O��N�%�����!�&�7�0Vbn!�3?IoF�ÙFë����"���
o_�� �V�D�8��OՄs�y�}�������	�sM?�d���}p(m���`�b��:J:�����`����ُwm_3�M~/��J�]W����i�h�&DҼ�B��0J��8K�5���P�9`�0�~���Jρ���+����^�x���k2q��.O�+�/�}7*�T�e�MZ��~M��#����Eg�Oq^��F�6�6�f@�M�NLC��U�6���M��w/3)�&�Eޓ8�۔�z�CzC��'��@�Gs��Lz����"m�`�kv�y|�n�Sc��-��Q��nC�Q�=��]s���EFS�j���B���?/����X$8J�`e�9^��[H�v��1}(]n����zw�� �yF����<f�C�Ǐ��~KZ�^�/ �j�dK[�zON`��?te�5�hT���m�X�@f�#�a����߉�jp��0r�
��e���������(0b�YrW]���L �'PUޡ��P�aa��y��?!1��w����u=�l�Ԋҫ޵�na�.�[�w�,��?��8P��.~%N����n���wѥ)����0�l�G��YR�:��ܤ��	P��N�[�+T�]W ʫ���M����C��(����cr_.�$w�
zq�HXg]`�>��Y%y5�t��~g34�"j(\{�k��	� ���q�!:��sфX̔�8iY�f��5�m�O���j^>X��	��tC����=s���,D�tF�ǣW�L�h��3�d�/��s�IN[S��#��_1pUڱ�T/G�l����	3�ʠ��X7Ht]�6a}�@�K����yn ��.�1�P`]���e
�<��gg%������EA����!�L�29��v?��y��1W�T+`fB����MՎ�EXZ�λ_���5`f���.Z�r(�A-V�����z�i��9t�n��c%)+�y��K_mk�Ǜ�fD�4����~�w��|�3�ב�܂}�Ҩ�A*�
o����~7�Zv��8Ԙ�'L���>ۈK�T��8C1g ��P �C>IN�i��e���0��s�`�|��#I;�e~���JR�na�?�I���X$O
`�(O#E�P�ͯG��N��QZU�b���5�=��+�}�+�[ݟ(7�>� ��-���."�F�2�f�yR�wW���9�Av��Kf���x4�ʟ��i%����_�!'��+�Lst��0��b��z���ԩ�۟���g8j��8
2���)���>��?*|��JR6/!k�҄&��^(�('�}�~O���m~z�&T���Z	0�/7���6Z
������s�!~�`=YC��F��#Z9�k���ID��`U��?����~i|b�A�YԮ�}�yr,[���Κ�-�����3{��~P���'�6�;^][tQ�$(�&K��CW|�HdyB/�C��m�|�k"�cY�9ɽ1<.��m�y$0;�D�"k����:.����B�ݮϋOF��>Sd�Mu�]��:����' ���:!�Xh�v����W�4C�БT�	�ð_�c�pB� �	'��@���Uu �vz�c"���-N��c���H�{Vā�"��8�zq9�W�����
��/��.�)E��m���Y�w���O:���o+_�~�K�O���DH�|7�۰X��<���"FyeMMv�r����-�r�Wah�2О�D���_"�~y4��_��:K�}����L��	�K���.D)�7l]Kz�v�m��Z)�^EK^~�:fe��8��/��6�J���%x���J���+0؈�b��:�f��_H�Qs�*�4�g�臄��I�uk�.f�F@F�H�)���36��qLN�wf����10u!�/dO�E�ߝ̂]��mx�!o�yMMAƎ/�[�$����5�ͩb�|�����L��"Mg��4���t�=�����ή�3�+�'����YF��"iе{����W?q��k
���x��d�n��wK�����4_w�A�{Q(HR�o������f'��@�J̗����+�س��Z�l��G���k�6��H렝^�6�_:=[G�rOO�BzV��e�gQo-}����>�s=m�	f�=�O�r�Ķ�yo�������tl��l����@s�4����?;�E��H(a;yp�`�s��$�'�* �nc{#D�d���U�Wcb�6�g�D
���4�������m��)
�ټ��KG2�����á-^.<B� P�3\ծ�+��[�Nu�3�|���wim��2�I�I��$�	����b�K����+7%�q�V|V�.�c̝��0ӿl	��y�6��|M��8�M�aOhR��jcZ�4RQ�H�0-�Ȏ!���0�iʺl2p`&��+ �~4V��j�ќr�t���T}I��#���M($����ҺIK�lڪ!c���O�­���O���K��svK^�W�9ᣨ���|�G�)T�q��Ȝ]�X����uK7���.#�Ҧ����R�0E[��:6��yY�֌�Ό�N y5��$O.��v@�����vV����Lk͠��۹b��W�O ��"zr�"n*tq�V����͒;���
l��]�L����؍�æM�.��g>��zɠS&��f�%j@멎F��N[�=y�z��䯥���ג����r��"�2�����1ƫ}.�F��r���s�bP���Llհ�eN�[��8B_��2���!�c_݋V��/y3ㄬO��Y*)J�
��Ԩ�������������-c�V$�
9��@{�:\d����F��3�ҙ���=52𯱽@��R��AUk&�ۄ�P���@،���!󎗨�~Dє�C`#����q;�%q�:�Vv���ɛ�HU�:ȅ+^z��y�"y��$��ֽ����䈤/4������)��,l{��j-��ڙ.Q����VF��Wх��� �ypE1|TvI�υ���ﶆ�5G��0 ���CV*�} #�.T��b4ߵ�%�c�a�O&A>4�^�=5��x��6SO��.J�D.�ZO(F����0��*�"�����*�)i�&���:$�Gþ�;��M�d8����Fm���Q�S��JnS{�o���[/Sj���u��h����,^���|���-���	��&^Kܑ��=u��!G��c=�NU{C�KoƔK���72� ��D�	�z��MvM���/^NZ9o��/&y��)m�ņ�x�vW�'��+S���׀B��_H.����P�4c��zY�����f���f�I�`(i$��@�D����j�A�Ar��+_�(���s�� gk�~�P��)�����ǥA;�u3a9p����J�˝�_���䤥�1M�ʒA�c�J�'�,0�
�f�̌z@1>Z�vN3t�� ���l���aO�9 �����>�ՄP�T�y��n�t�`T�����UI"�^>�h�>E���tޮ�p	J�s�4}6�@;��x��#[7�nx����-Cq�_�߿}���USg5��ձ��H|F@з)�2���|)��C>1^�$���yz�7�k��Qc�Y��F��X�`�[ 넻{�_��d�dC��%UQQb�j�]�B�5�`S���UW��4P&4��������/������%2ߚq='�>i�7�A�#M��C���wn{2W��u�.�9KM�+��Gc��(�7-O�ڣ`�v����@kfDG v���Z���Y�/��D������2Y�;�&���b�hk�3N�\���Y��x6��5���'�V�'��uz��d:H1_D<p���?MA�"L�cx@����	�6�!���非&^A���o��2G���*��;�b�F�Ĭb�t��e��Ts�2l�؂��9e�)L��dí?G\2�>�������q���XL�~ά�S��]b����;7K*��q�hT�w��JvM��d��|�K�gƲ9����R�EM� sjJ��x�/]���q�gKrRS��{0�t_������e�Y���:u]C��{���<_o��\�k�mKJ^��l������ tRi��.-�
�����$�K �c�
�V�W�h��kr`��L��T��VOv�+�r�Eܨ[u^���%��~j;����N��E1w5�����bR�5[�D�1��
���s��yJ]#��2&�,��\q7�>=�=o���s�"rL�?�Q�����z���1P=l�d��e&��*A�q��;C/��1R����Uϻ���W{�*R޷5��v�T���v��&� ���nd�C�[�J�����\�v�i��Yk�������qb��t�v��2
<����˪�Fn��l�y�X��\mml�i�$��Z�C�In�N���rI��ԟV�
���:C��j�.������Q�� ����:(ސ�� �e>?7k�Sݲ��Nb�fv*G%��W��O������bo�<�z�>�|��8����y� �D꽌�A#OX���g��h���gA7�0�
�h2�*ռ;,<��Y`���O=�-Q�x��H�e� O_���+~m�o�6�)kG,~���E�&�w�Q{�`ߢ'�
���^_9#QD�q�B� u����7�3Kx���}�Sʠ`-$'���ަ�e���ؚ��M^��p��ݲ��!ǟ_� |��mI��w#�(����P�W�Ycr���9�`�a2������['�&{2c�)�Cam=�u�4�§�0�s"u[��
�Y�s����x2���L=�)U{0G7��B�E,A�i����B}���t�c���w,�9����@��\8��$�8����FסU�5�/Π��o8����, ��6�|�˓ �i�U~���'F@	�*3��!����嗶zJ�$�����T
�_b���P��b�������C���dH-�J)�����;kI���+��κs����������~w(�l���Nn���@�Z�g���}˶����!��+/t%��cOl]6\j�^�@�Cs��z�G_3+������2rn�	괍1�7�2�Z�`Ş:W�_�'�Ȓm����{W<?������t_
���QA3��QS3ą�~m��eB��G�{2���3�ק�&o�u��5��p�g���� �%���H��T���v�Y���^3d�^[��Lg����<�ԆwBFd���Pq���\�ʒCˁYoy�	��V|��"I����(�3:h�jyo�Y%����M%J��M��Q-Q!�j�!�aJ�=��WS��x�o����y�>�YҨ���R�T7��$���9����ۤZzG��@I�r�[-TM�2Ks�����d:����Ǫ	A#���ئ��.��2�t�܁�ސ��
v��4��14�H�}�x������}`]B�����!���#��[̪z6���<mxxx�uLH���ܔ�Tq�w`FO22F"�R��v�?�ʟ
��#ť83L���:��2�HY�Y�K�1Fvx=!�{���f r��J҈��.2�A˶�k�9z��W C"E��!5��#�<mz��p� ?��;�����2K8T��T�]��^�Q���_����!����[=F���i5��'�����M��BuT�:�z�����-����[��-3���j�vq]ٸ��/;A	x�,򺵤*?���SL9w�W�L�l�%�U���_+A�C�IP�Tjk����*���{��ZDk���|�pĮw��˯Y�Dl
M}!�#�5�ٯV"ri�Wt�x�����{�D���p�HM� ��+���ޭC�0<c�r9d��^^~"i�?���I'{���w\_����+>mk>����eU��!e�01��m?��̶F����o!3�%�T��˼A���)܈xp5��gp��~	�eq�0����V������;Ts�Ǟz �9*�M��u����hS|~��v�
O������k�c�j�ؖ��hF�;*����v�슝���#���,O���-%�%�`]�������k�ý�v6��WGǻq=�'J9p��"*q1��j"��eg˚��gw<�Ĳ��|�&9���� ߝ���������>����ܻ*�_�|���)�O
����;���e;P��6V͹=�4*;���o�<�`3P��J��gC/@�P�Y���nhe�m����X�[�"�liU_�ns`�F�c[+O]��^ ��O9M��hϏ��i��`����sH�R
N[,k�=k����v�۩�,!�$�-���TY��џ��B��8m�cG�.e۵ak���_�����Cj\R=����9���zO���r(�Y������a`Ƞ�����a��VX|��:���+\�b�к�,E�mnz$�+$�p����t�ssu�RFҝ�]��~'D��\o�er��P�QN��#�Kt��������>�%b��Bh7�S�꒕j�r�H��4�Vrua@ϑ���jcN&�]CE��khl��6�j${z�6t$�W6����+�������to��ϔ���I$~\#�QA���/����z��\��Z�n 
��]�#/�h�g"q?���F����廤�8��\��`5���9㏀V_�gV�x��|����k*ҩT�8ao/Ij#�:D����
�z]<Vw�/8w,v�b$%�n�ԝFΞ����Qe�4�]��Xj�9-�1�_�$v^��� n9�x%a��x(=uZ�������+�b�R����..Zz�7V��Q�PP��Cs�c�͐Sv)s�r_%57!���B����R�W��a'�2`A��b�7T��"q�����	�H�	p�/{�i�E��X
�4�ÙsQ�뷐"G�%�5��O~k��_��C-��J�� F~k.�au�)�Y���2�DG,�N@�:D�!b&QQ�h�m�OQ~��y+�IW8+� 2gFG0��N.�#q��c��pC����.`���Hy�m�!���A���r������j���a�_�����Il�aϰt�����볺F>�)(�ԟ%X\cwH&L w�ߨ�E(+X����<��������Z��V�gI��lZ
�G(�Nգ=�S1{f�j[&N-~���""���GCu'�ؾؑ���l����F��R�yq�V���1�z��vԫjΫ�-}D���@�M$����mY��v���5D�@���L3����w>lNj����6��g]��?�pY��P����Dq2�<�Ĩ){�΅Xρ}(��e�V�����m����ߠ����0j����@[���
G�5E�&U���0�m,��žV%�C(���)ߜ?S�p��^��_g�ثL$AO
� ]]��$w���6��ds���v�;��3d�1*������ݲv�d�[���j8.�1I��}�eN�n-�_g�b��~���rl!<xGB�J��gB�7�"�`#~{VÍ�ֶ{;� <��`o���T[h�E��X���}�����~6u-��asf0b�;���9(�A64l��,�������'B3�e��N�O~��ZV� �o]$e#��T���#d��Y�|@��=��$���b9� �wv��-:=�L����Q��)�'V	A��hX2d�D�AQ��[�L�\�G]��	�4ѩ�M�DǬ��׭���R�9�89�;k��}��,�ę�.Y\Fɻ��":��@�{Z;]²L�u_[�g�/��ٍx@:��e������3�E9�Eߺ��w�& ɡBA���q8���Qt���I���(۰x��]z�|i܄T5��>�C��~qB�Ӟ8�%+\"��%�^�n}�L�cp�on�qM��z�t,[��]T�(򵙯�7xϳ�d�~+x���@��*�ﱇ'ΪX�b��{�e�7.N5V�61=i4��	)wCT��.�C\����Cׅv�O��������tZvj���=8�)pQiW~v�����Gۂ�<Stn .`5='i��(����, ��t����mZR��(������b�E����̶�3�"Ì78�)�_nV�(��5�)--�f�=���(~�_�����8ey���z�[�*{(%��숾.z��j���6ZӇ�
�3x�{Q/-dje [l�P��a�yL�
�������.���ӽ���_���|��k9��T�� �:��ym4�5yG�24��r[%�@tA��vR�X��;��}�O(x��}y��j�瞪�
�v4O�KN�s��VW�f7*�vo�@.3�`�<����J]��y"��75�OV�E����=��<$^O����)q2�t8��b�Ci=�9�z������#�c¯掆�mzb�|�?�c=W�����i�#�������LX���m���'(qRl7��63P���F֒��g;�hb��h���wx~
��DIͻ�_�l�b�-�LD(ߦ4lyU���,��4:�����I�r��4ଋ��7+b���jI��J��2C?��zm����0uGx��cZ�[�G���)����� ҟ�ZĚ�a��{��P��
L���
W���PJ\"��;!eB.Xu�5M��]E���%h���,g���s�<z[�����$����iFC+��l�{�����r h����~���e�>9�Y�<)(��(�)/F�s���D��r^�X�d@mn�u>g��:�q!�<��գ���u�̓`���XG�J�>��uV3w.�/�zw���?`�G������@V�?DO)��A&�Ì$��H:�M٭=*f��(��9 C��f���Jt)G�r��[L����F�Ll;�}�E�]T�-�N��I��PA�h�9�����05���ۉP�� e-4��t�j��D%��p	��N:��g�`��O���,��9�J��i���|V�.�c9�Ƌ���>��#�u$���Jl���t�`�J_|��4I%�pfT���0~i��ʈB��x4��e�}�ߘ�1OC���qȰ�pY*�8s�+|����x�kB��)@:8h�H�L7$�2vH�t�����������ͱ��@fU�t�:Bz�=�j�g������2�ۖ�r���k�vfۍ)&�U�=�R!q�{Ȍ�ei���l�Fc��}i�����oh�$0�"�? �
��0�l,��+�����#j����,����fKM��E��Y��>>�ʌ��}	��y7�bi���D�iz�a�`�?�>��s�-K2��@�ﺦ��-��9�zE'dɁ(�|�}��`��|�[��u+|���Б��^�M�~��������6���de%�5>�T�(([���Z�l�G�:���,%hw�c�N� wKw��M(h8k)/F��݈T����z<Fb������H��y)OV�x�<��|=���/�dw%��7����K92��.�<��L�Hţc�T!��y�OHM<HSK`F/���"��e����p@���m��$��x1�A�g��  �n�:�O���M����{�����|�0A��ɧrucW��˦[�����Jɷ�z��� )��nz��|��`$�>��r���QZ=&o�����e�>��:�2�X���83��ftw� m�ˇ��b��y��_N��{!�!����0TC$@���GO�Tw�
��@��$����;�\"@��̂%0i��g�J�4��.�=�;�fan<8)=�svʘ�6���gW�!m���g&��(~RN�
Z߁�D'L��������0��g[y?�)3������r3�R�:��`��}�!W�d`�"5A�=Hg��l�)@�mL�Hv�Z[�O8���?,�Lp�|��+%T+Y�:�6;{�Vi
&C�6xƾ=��J6�|����L/�W X͝�J*��{��N1�l��!i���*~ *��i��(�����ϭm���"��}̴%��z�4<F��'��
���z�Y��'r�לe7��@�eZ/"���_��"���E�l����C~�]�m�c��"�n��w��$�φ�A]��O�A�c�@��Ą��0��͉|8�X�m�v�lvQ�����^C�g��ny�v��Z$E�o�߂%eo����\z�e�aS'��|���8aH<V���Z+�jd�W��]*�$	�E��j�����Q3����$�)�Ν 
<����k�]��
�1�Oh!vg�`�J!>�6l �\z�$�d��w9S�/'K}ٍ$���#9����聖(��gv�0����Q�Ad�pR�/�@�tG�����s����'�JM�jo!-�5�ۡ8�Vܶ��f���k������ �*�|���.�p�U��o:dϷl��T���o0�6Ҷ�Zb����Ba�=�*t�"u^1��p귁,Mؽ�D.��<���ϗ�mrk����ҔcIu��LP�oy/�T�K�rb����hBI�� H��{,g[m����:��1{�-�p��,΅�ej�>�E$��k*a��n����>��v�'VV�`���d��ލ'8L��.�G�MH������S�]���Uguʻ8G�i
/���Mٝ�*-�����K����ͧ�wK��N����X2���4'����n��@Hc�q+���5�h�_�wyP2_~v�hb��*���Q�[ybJ�	�TX����������(X^�4KȺ����F�15�g1n�=kX��Z]��V8�zҹ�;g���
�=�v�4�~J_���@&��������۽=h�֛Y��hP��.[�! �Ԣ��q�U[����7K�5����,c�m��_�1���'��a�`usoCZ�%���&�2�@�>�DѮ.�m?��,�B�S?���o�MZ0�!�1�ɐwE����lg\����4z���h��-{���SY��%�~��&#����&����^mB!Osp}���٣-�F��a�薻��o�Az���z��pwሑ�1~t�^�j����7�3�,ֳ�TF��St�7�2�>v�y����gf���X�U�G�(�كu��/@������$}�lL����K�����H���{c�f.�~-]w�ɧHE��,C�4ӊ��G}����32�ݣJd���)q�㺢����ø�=HS��b�zG�5DMuî�=Q�Y� ������N�Y���k m����z�`І�/��D�?f(�.w�W��h'�1�Q���Y�A�FNԉ�: _�cc�ڒ��&wP�M���xR6�5�3��L*���A�`W)3�	U��r1�6E���r�R�EUd�{B�4@��<%gJ{WA���%��B0
̡���);?CS�j���k�d]�rA������  x��Pd�AJ�̹3��*���ǲy%��Ԯ`�����J�uW�k ��8�� ����Ď+J��9[tN�{�  3�4��W�J��x�K�����h��ʛs8���u����a�;�ϲ�� ���3֮>���s�ИaLp��jY]���7kխvd���-���<&?���|k\HF�=F@�Σ�N&�	w���B�9u�m��h����'�bp���jإ2�h�_<g�M��Yz�v� �e���m�ͪw�%�'��;]w!zW�,Ad��͖��*��
�_Q�>+B��\��V]Ɩ '=y[�Bq7�.w;dT4gU�s��+Ї�P7�0�Z�V�"�D`��r�&�n��pLXL���WEfM�z*=�XKհ/?��T&��V?�;E8�b9��2���@�`˚#�tl��Pj�����N`��k��4��^��+F `��5x�9G���@:���	�v�#�����I�a�/��sP<I�I�ʈ�u�Ko�e%A���w���Vg�Qz�����dsh��J���,�Ifo_F1�?����O����d~V�ف=F=��k���e���Ns�k4��zĆ]~��#g{����[��%�%��*j�7�y��*t̺	x\tȡf,��g�/�c�uSSzT��<x��&#x8�&��<F�9� �*XZ�,�;�t��Aħα�/h���\��z�JQl�x�^�}B�lb������{���EnZ9x���Of�WJP*F�6���
�^�v.T|?XH����_h��R����,��iD����HY�bNb�A�>
? 7�x�zi0A����3����)`�2 F��r��Mt�x���T~�#��t���OVA�%U�CPf�Ģaqi����C��mޔ^*��y�.]Y��>�[������]��G���l��S�O���\���v��Q�`�82Y�<�f�W��[� �*��FY����?�s����o��,����xP�<�x���6Y�NOd����g������4���'�uĸ"^��q`WgE���푣b����F��)&��@��/8�؋}��E��\MH]�GuT�!.�q��q��Υ�}y�L+OQ����o�ٻϋ��
S ��,e��8!���	������_��+4$�X_\�<O\��"�=[�B�N��?���(����-�;��u�CSz#z\5�w`��:0z�g���,\�^��/�[H!��t7�.�>-�j2����*��_��i��*�#'C8F��B�bs����.C��sUJ����MS"�Ǘ��&�I��O�4%^����@D�P�r�����O�wl��ڊ�x�2&�]ߢ�YI|�����j��G�ӓX�P�V���-ha8�δ����*������E��>��1�*���U��p8�4A�hL�4�Ӽ�WQ��i�BP�}�rr�7� ��.�'�6N	+� _��-�ս�UЎ�c�� c��نQ�!i5JW	'%��ig8�����jC��r�^��k[�L�����CX�S2u�����L�)��q�r@*L,W�0_@ eɚ&`jPFE����>ao|C>��q3N�[yl����eݟ��3���v�nfJ&�JY����$��v����u_7�����5��5�q�Ɗn�s(
�a u�������=g7����Dn�N���n���+v�@97�F��H���j�#'֌���);�P�]ݧ���R�W�/s�50͆nrY�-tM��6]����6I�5�n2�x����}D������5n������tF��/N l�Z"���#����K�rm���̦���a}�����dk��۷��J�k����vCM���[�������	!���/4q�������t��4�i�q�,�&p���0�����b%��K�r�.�`9QA!\�@߲N�T�6��&f��#��+A��"يԈ��-~���f6֓[7�uC���7����~�{Xkm�z��!�y�]i��T�p��N�ɸ>PC�����FzKO��'H5}���,M��w3>��¡�*1L�(o��R�%��� R��?td(:	p�_㽠RK���'N2cA7A7d�;��˧-K�Z�h�2+J�2��'�;�W彧������'����u�HD������Cr�Y '��P9�W�\3�2߭H����{��MJŢSF�{��J�������6�N�������_7yƕ���m;�j>���k��k~�Y9G�v[����sg n�|s� �w��u��R?�/��1�']m����W.0�\nH#Zr����r�(���qY��W��T�p���t��IH�a��Q8}K�K��Nh�,���6�P�<�t���}6\Py�A��v�#�k�U`hd��>d�Ѐg�&��M��)\l��	�=7��������v�*��D�pW��m��+���?O�zYW�z���/ׇ@����o���`����%%��Vے��
�ҥ`����Mcb�Z.RŸ�M��{�/���0���fl�^�d���񆠏T�6cÀ4/���i��-����oF!����]6X���m�BC�y��cwS;iK�6ni�JI�Ap�����"�$�Y�Hkƶ�n-,2I������e�o"%�m�d<h�5C'�7f�+����!O�|$G���p�z@��R���kl�r/�L��s�!��)s���_������,X�Rb��L�׀(v�LHL	GW��fjK�`��/�;��(�$φ:�)�`��2uI0���D��Z�̅��'7�[�4��tٻ���؉}E��dd`�r��J�W����M_�Z�o���J-T#wu�����@���3Dc<@gP�0F���]���F����?�^�H>ͻ�+ߤ��h�^ L�(���/̞cQ������zsu� �Ʊ_��;�0(4gf�XV�Y�f�C�}���S`Vh�f1E��-"jO(;���H��\U��<��9{��@ ������Lb���lBK3:�o,�~�x
��w�uaJ!ż�xۃS�3s�����h N�0x��RGA#�X��6�|���G��~���7?q���ij�+\���*��K�5�7���̽��H�r��<8��㭈F���f���O}_��5	��6P�����#�H�|t�HU�B-��9kh��nd��&o�C�6y=V�[�.<�sEa��B�Qp�*"@�^���x�D�$��unLҽ���C�F���gw��&�(��4���u���ɱ��(��tj�l���/���*�I�>�.W\�yO��:�r����[p�K[���P΁��	�UK(疁A Ǉ]ճ����屽lE�����Ÿ1h�+Rv��W��86&��9�l (u3���|���6"�������-�c�Fl�|��HOFݓ����&�H$���;���o~���u�-[��dn�R9
xf뎆\��{-���Q�(�����H�ʤ:�'��9 ,������Ųb']�p�a����V�5�ן�)�����p$q[@�������)�g��ӌ}J|�d��4y�y�#\��̐ �!3JOND�v: Zp���O �#��;�6��Y��A��O��C�-�8�Esni��cq������E5���~n����Nl�΅�y*����!�Ő�-��뗳�e�|�e��ӟ$�!a��T셣)�
������2�ǃ�q�*�.k��Y^U�Z@��s=���vk~�Ts�17����`��
���$����8�=x~E|L��,������6���E0�z"�st�����z�	�0�5�%�G���<0�asap�`
Z��^�Q7�d�3�y��ܠ�����s����}�>RAC����0=�@���C�͞���sH���~��e\����5�-�fNg�Fms;*��lB����2�^�\���
@HJ����o[¬�L���F���G�G��j��!���R����t� u�r���ž��*��do�'�10�q�����b��5�?����>M����W�XI�iQ/5p7�V8z�*L����	�z�X"�COt5����c����%�1���_���1(�O��N�w暀��>��0m9ZQ�e6�%�8�:zyY�{k�iPP����ٽ\a��+/�zW9R5�4-�B�ÌT�웋���\l��rSB��N�/��&}e�P*YH�j1��*#���B�|�x;��khv~ü���qK�+�>��0`XC�������D����vXY| �7=T�s���dfF��ё���쉵rQ|�CX����)*���Q�<���Î���7sJ�4��\4"t���C+QiA�a`��`�0�9>��'}W�P�9si_��bz�|d����oT�>��L-k_�Е���9!��ܢ�;�I��_����`M�J�w*����@��E�{�<�[���}�;$�ɆƟ��xǉ{b8�����x`?n�v�P��Y�dg���?�e���ɤ��p��ۅN6}��W�Qb7:�6R���OV����+�r�,J�澮x��@��Sg��o�is:Qu���� /c��UB?3����Z.7H�6��:#��"͕��� ^�	�]��WY���yMgi:qؚ3�7}"o_Id���0) ո/��NhL�L��?3rW�u�O�m*�l��\�~�9�7�I65���ʪٺ"�1�F&^�8-�+f�`���:MWkwFFA���*��tp�2/AA�!
Hg�e�.1ښ ��Tj��\K��sʩwW���p=ɚ�? }N�����⎭!r��F�$�Mc ��6�'T�Ț��X.:��3H� 1���e��G5����������'�{�ՅsZ���988�-��n�/��I�ָ������k�����&�W��g�0Nb���tC�Ȱ!�/_a��iT��w�[Jc��|/�N$�W���l��<q�'0n�=��lWFg�\��B��JD��u]��>}zo�Q|"ݕO)��5[��k˺ײ�z�,7�l��f���L�`�\��ZU���o-��0D,<sl�k�K���^dz}|���O�È�}�?��G\���`��4)\�j^i��\E�����Qiđ��nvSj�$�zy{RY��bӇ�3#��H<-h���-�i\�$��d����8��)�����l�jWRƻ.]�[,-6�E�:Aj*��V�XB')+�|�+>I�P�+������J�F�ɞ�a��̎��_�����\���օlw���"��x�@(yYs;�G�+���.�^y���[�n�t?���ߢ@��G	V�}։+�b��Q�;!	���4E���(�16_xU��E�Jqi����25;��^�4o�'�V�w�Frcͼ���M�,Qlx��'�i���u�����(W�=�k�8F�>xs��=G�K����o���(H���Gp��r܎�]��B��ea�V�����4�x5)bC�&t���UV����X��44�1S�m��a��H��4���I��|�|����r��g�zU�(x�Z��(�=��d٣H�h��l�)W�lj���-K�6�|m�_��*ܵ����T�⽺��p�^�[���3#Y���9��;�Q�ä�e������M+�Iˇ�(��<`Q�/*
�,׵���h�z=fE����*�&��<�|��,-A�<�嫁Y�`����@Tg�C�t�F9l��+z�#����N�#\���f1�զNb�"J`��e�I9�i�Z�u3g!���~t�S�0�f�L��fO���G�Y��{bN`��.��#��_{�Ԗ�m7et�
�/\M��8�_ȎZJt��r��R��r��/qNo�v�C
@R��� 6|�<�Kj�%�ƃ"9gH��0�"�E���"���󓩵�x5�|��{��b��n�e9�Q�^�K�7����uQ�v����^I��j����1�B��Qf��"�T�%D�!� 0�Ѭ��C���|��/^��/�t5�S+���~5�ס�x
r�W����1�}����į�r7P�+� ػ|����!:�DyZ@wa����Inے���ֶn��?���k����n���}�~��\�v+")������L0ٕר�/�{C��=����=/����|X��T������X!�]�3]C'��0���B4E����q��RI���T�U�.�d�D�\Ì����/A�F�0G�co]!t.Y2�.[9J;8�$7.i۰��O�����9��B�u�}�h5lN� �d��;
ߔ;�~�����1��bql�hi�+jX^��n3�)�i�9�A�E�[��d����Ubmб�6-��,�>C܅��Yn�_7c\t`��s�v权�	�5D%X���f���6;x��l\�� �A���AP�y��O��qI�&�ݯ[�V(��P�$�Ч�ب_&s`7�1	�����}.�ȆF[9t&m�s����Q��= N�#D��Ҙ���Ň�Lq� :�&�j���Y�9�-��� �:�
S S=gϛ�D�,��Q{q��{��n�e��"���G��u�^�o�NC�J�*���3R�<�٣�����_��4�Ťa4�[������� 'U_#pQ���q�2�=�mQr%���;�m� �uvXQ�@���4��S��&l~��3�����";����}Xj~e�\�	�u�(�CU� X��1T���J3e�]A1�/�����~��nX�;�L�ˡ Π��m={�p{f���5�w�X1�^����˴�N)��T�A&N��v�XJ=�%.�|#.u�g�U	�ї��7�8)�/P�9�ӹ�s;kޱ�Q+u�G���/VQI
y�BU�}S�ܭt�����h��|�@԰i��\� ��S���}�٠�t�^̋&��7X?tdNY7`�P	E���>0S��HS$���kcp�GԠ{8ƥZ ��#�	C������q�׆���A)�w�V`�k�����9��1����{Ǘ��m���(��搝-px�9<H��G~�zOҕf��A�QlA�� �D{�M+��CO�-��!84��h������@�7D�Y^��Z/7�Mp	�lE�^���~�$Z�H��9Qv����bm���/b'�p���7�dh���4F����=; ^���ˇ!_s�V!��6�2 g&��,K�;-���g�uV��Cf^�Ў�"5�w����ͤC~]{�9!G���x��yD�#BЭW��1��ٝ�bS�����j��ǜǱ?��XM��8El���t��ιNՑ����v��p*�w���k�G�S��Hm�Tͦ	���'��F��UO�'�Cin�?�(�#�He�~�ӧ��=q��b�*����4t��v����v	YR�-yu}��J)O�╅�6[�n��^�	���/����ZDЍ���:��8��rM�{9����-������%`�&�4���N"�uB���UԘ�%Nr,��R�(-��k�n[	���]�{2B{�{��EdrXC����sY;E#��_��G�Z����ł?|���!G���b��
��"ń��GT8��F���2ፉ�~5���� �{�@�*{sI��0��ʴ b��g̪��\a0�͌��8�>�٣" g2i�Ț��T�\݈��z�":��yY!��<�rg{N�fu�h��Av5�J�[6I�rr��;���*��
�[�w��@��`����p<o��|��)���L�;3�d�yY���f�d�V_�ޅq�#�(���2S�����:墪��^`m�1�}XJW�n�X�Y�C�w����,�	�E�8O��n��A=�rH�n�_=3�=���?윥��A-��ɤ�.ȐRӻ��%�,���OS:?��2]-W�U~r��`I�Ns�x@>J^8-�����D�)<��ٝ�~�5���g�"����Â�g^�r�fK$t��pHI$��#:���@|:X�+/��r3���Dϸܟ'���$� ��cz<��W`���h{LwACa�,>^\W����6�ô�[b�r�{47�^J/x�gtA8�7�5"��]]RJlIH	\�	D=���������� 7��Wթ��i	1���sO�|���N�q����*[X;������D7L��X��:�1��n�2��ь@$K&��A���m�D��*�O���K!J���;�Ǿ4�E8��N��Ҟk�|eFs`'+���Zr_��-t��xHE*#���(��C`��Njة�� �BNJ��x���(�µ�xV�=y%v<�r3���l�Z��	������ :�^��d���[NA���|�����C�ҹ�h�-#XK��ZoT���C��_3b���`D��bh�蜐ڼ4��o�*>�,�6�2|l�(,Z`�l��d�6�<�w5x�lJ�sW�J�Pc�T7Yٲ��7&V�u�)�p9��U�]�k[�]6���2>3�!é��C<d����GO���	@R�_��óŭ���T�@`RT4����	����s~�E���
�y7�m+��M���<G�J+"�P���Ej�K��wf���0�\���|e����376}@�u,I����b��Cv���.xvJ=�دt�I��"�q�E�_.�RKAJ����@��'0��\���Y-��G�x�����s?�N�}\����g w��{/��<oTEI�I3�(պ��;�����L����þ��[O�R.��e�6�8���p;�e��N��(�%���T¥PY�����qA�[{��	I~a���ib��NM
�����-��t]uh��{%�"Գ5�cy0$;t�SLf����u���Q��4c���<ި+��aL�CK��$ga����h�>��~���nv�oF⥃W|!N���p��XwvS;���X�f$i����O9�aCEy�l� ����T���n7���8=2nThB�pZB���ϣ�aY�?��j�&8|{{Bh5�[SH��D��1p����u%�*��,�<��:]�|ل�BQ�);��z�4��s���n��Ha��+6I��|���Y��c��l��V{Ʈ�	����
��\?�v��]tpі	֬����~�	�d�(�{�S%����:LA���a�3�'���.��dn�dD���k�p�ړG^y�7p�d9��=�+��V�����X|�v�P"c��R��l�'��X�1P�@<lyaSB2r���a3��v��gVD����ֶ�dD��[(��k��鐎�����H�ҘwJ�k]�A�><����e�鲟� @tJT����gC���.��"�~?�16�5z���S�����,H"�T��4�Ҧ�s宒�Z��T�/{�DZ�CP��`33MJlA}��J��P��a�3�
@5�	�oZ�IE���Z�u
��Lp�M�4P��t3�Uc���z�m��Xӄ+Ȑ׫�F!at�d��J���i ��I���JWpN^�)z+m4��{/g�8AC�9�ȅG�x��/\,�*��7�-�,��9x�h&@co���js+
&����z-�1.8Q����k仕<%/�C�>�p�e���"��qJ��K�}k�u;\�ˠ|eO$̮�ߦ]��k'gPg
��P�F��,��q�"�%EEy�C?��7�Q�8K����m�QT��L�������8
�|J(}�L�#&����/ db�R�nc�f���.��Nn%��b(:�ܧ���a>��x՟+��'��� TX4�^kO�a�գ��%�_�А�2��,*���-�j	�ڡ����8�dd;���vn�X��|c	,ri4���JfMq6�bh6��z��AC�5�5��[�7#��� K����`��Tn��`�-�.�i�,�u����u8�����3�5G��\�9{`���N�s��u��H�ZU�
�Ŵ'�
h=���s$09b�y��V����3}H/e��b�&!�x���@iBw���/,j���k�4ӈ���5��^G}�8�]��n���?�۸|�C��ӕӸ>� �D��Vu�L|�b��A�[��,��T�G�����/5 �p�d�;'Ѫo�֖��w�)��/|0>����������y�\��)����+�&0+�D5�_OK ��w����u�B$`���=]'��~X�y�։�S��a2_�t������2J���C��E�P�ESjY�/��������LOn�ծE����%$<�{���l�.��p ���?ez	
)��B����P8f��ܤ�1xc�#�&qRWb�A��������J�S5�^ u�uC�kc��ii|19o�)^��YB���~{}�{>޿�1W��p����wK>P(�;d�Pv
�Á��	��{����Y�\|'�x�%���e����M�p�#�'�!�R�ѻ�:���v���v4S'�
��	3o1C9��bc�q�ƿEݿȧ��k��v� I|�_��+��qf�'�ZB�ӵ��춵���׶�v��yF �bU0�-�#�_��\`�@Q<��|Ұ��J�Ǐ��H06o��7�u�!��L��Y�'�a�;��IP���--ng9Ӫ�r�������_������\���|��9ĥ0���HK���$_�����dh��K{U-�ew��u�8��#��of��ʘ�/�y�"~�x�7�j%Q2���
9������^�ϵ��u�zx�������;�7�$�t�On�I!i��oM*/��@��^}��g��!sӷ��a�����p�r�=��KaǊ�~����n�T
{.(� �&�~+���+��r���p�(�(%��qMK���m���	��/U��̍��4Nc�p^��K��1P�=�x���&tAd�V��G `*����kԙ�ݽC^c�a��f�jA�Wp��oI ��K���\�5����pv�Z��&��0�s�Κtb��?dV������;��C�%������e	[�Ll~�V�U�2S W�v�kZ?0@��Ym���5Z�V�+2�r��6�_Ǿ!W"�4��񵠀�=y _Ů ��.3�^�`�h�g97Ye�N��آ#����v��	lw?F�]I�bH����#ԧ�P>q�)�D�v댩a y�TS�髬�g�Lvu\Za�RK�-Z�~�=�an#��.C������j1��.v&Zɷ_���Ba����%�x������&��;z�t�ɹ�� Gc�"�)�p%jū��!7�t"�� >}mb��lp���;�3UlbYQN9�HTg�*G�k���q��	w ���(��q��D�c��R�Z�p��s����frC� C�D`�Q��ۓRj�w�w����m�VW�{+�*Ns��J{4b��'���L���r�ݼ�c(�D_7�)\j&��$�K�=�8�8���|x���zh!��,C��Q�m�6��� ��An��QD���j>��ϣ[�R�O�UI�~28�bۣ��Z0���J�0vL�E�Z��f�É��zJ�l���(Rl��9�P_�	���'%.x��)"ͼcu�O�<� �����oP�W�g������f���-�c���8��-D�9��O��\�I��h��Y�9�p���YO����WJ�l��v��/�S����t�Ԉ��΃M.�X��AQrs%����G���u���=���2�E謣� ��,Y�����������n����A������_���ծ��0T��Kh�
���J	�s��ρ����dO���L����#:-�E=
�ӓ?�po�?Ό���b��u�2\��FdC� A��O@�{����8�v��l��-�<+��,߼�^a9w�ky�*�U�j��5�}Z��3�4E�E(a��"[� Hj���lC�u�,.|#ԈD��{���pj7H{y*Z�P�^�f��� K��}�e.@�K�.dݎ���[y�5KF����q�I�'J������c�-l��{q�b$X�El_��|4�5~�q�W�����H�2ض^��H��M:
��PvW����g�s�,]��+������pg��l}�9��2l��9�H�#I�A���Vm���p77�<wXE�K���9;�j!�����
�����2�T	=tjF
D�U�s8{��,I��͖��h�t��}XP��)Rj�V6To���MËN��Ø�p���Y�W��M�U먏��k�dl�T�ɴD����VFEe��t��M*��g|�A�9JwN����.������!����{,TK����o? �Վ���j�S4�|��c^�5�k7���E`wX�؇���L�������Wc�:��f�,&�3���Eb�������i=� 5f����W,�l�)jA���g
b(�CϺ'�'��	]�Q� ��K?��{��j79�V�y�;QW��l"��
2��	w��46zz9n��<�[��m���|�V�"����u��n�3�p#��vn�Y>'PK͢hC���?CG����N�ʤ�1`�PرF���gX۵*a�"��_euTJ?�~~���e�Y���(�n�F��Vd�K)�f�A�a�������q��C|�b��g���[�q��Zf��?��H>�d��Ͳ�4vդ�]~�3e���o�6M(=���J�A�*��#�f������0[CN#�	�ϳheT�K�lrJ^�/ Lܿ��OcQ5ͅ��SDG���[�jPH��fA�+�5_��[δC~~��>iP���K��*G������ML3k�4��YLF-Z�7����:��[�{4�~:U��0!�� �ZV�1�U �_ғK�ܖ�m�%�A�V�{��
����8��a�D�AEڌ�'�oJ���mrT/u���!K���N�����k�<.�}N�ܪ��R�><��0������I��Y��k�	HC�V�(f�Fd�x�5b���%��1S����ܔ.m4����u�^L��A��ڻ8Ы�����B[��s5H�g�ޫ���,�@ H��g@��wK[E �ֱ���F�1�T`�O L�}7aП9WL���|�]s�L͏���%`��+R,�X�6-E�ݡR���└>��#�-̲�Fgʢ�9P�)`:Yl��22Y�n|T��w{D��U��e�I��SФs����{����?�%L?t�h}ni�'jm�DkKȑ��8$¸s��a��(\�L5	M�H�eG�IS�)�x�;�XA<v{��!|�i�=FeBJ�M��`��C'�zu[ ��!��^�lhp$�ʌ�~�,E�c#���`Gje�l��!>}8jZ)C6dY�H�o��L�f�������7�v��Ꝩ����0�i=؝u�|K�$!�4g�Y:+�}D����c|Ŧ�(�DY6���F�lf
�6g^�����=� �@j�ů�D��\�T*�f���T|����`^�,h�2@�޻��h�{BU�(cv�tb�4��!�YZ�m���oSh�5_�d�i����+G(���%��
rk���V����pܼ�U$���ה�F�o��!�RXp>�=.?<8�����D�C�?�%�}�'���$�����cտ���O9�	�ӧ�I�W ��Jc�+���=Y��v��a��Bܒ��##oF�+�-�^�*���a�Ƚ��YW$���֤2�ǜ9=~��:������2	��p�Nh���]!8��]�����W\��=͌���!1ؿ�^,�����`���]e��#3Œ�t�&���v	ݪ�M_�R�y��eR's�Ks�'��������*F��W:����h��.g\�]�%kK��#S
}�$MV�S�����!��51Oc��Fo�̄���+�?�r��oOh}�ITS�u	e�9Z�4gV;�/E�@��� �s�s��Уh�����⭸�|��
ks��\Q���źl(䋂#��@l��״� Q��~��O�-q�p =#8]~��z7/�h��vL�汌	�`�	腱���3`,#S�=�)�u�f��vu�U��m���i��+��7g�L���M�҇�5�r� ��8���q�����+;S�!Dh[R:�A�������ѥ���m�����]jA%'3>������t�IX&�1VORX��&>C��J���`a���b�siʖ���(�I$�3��EV�L�BBrud	�n���{m�F�^�j�I�z�Il���ȳ���E�{ڐ~��ߟ�>vS:�7`����J�֖BR���=�0����ٌ��nE[�A��,4��z�<T�z�� �Iuf�qY�'y��`x�,2+�Բ�D���:��p��FCN>� Tߣ���D��)��Y�c.��{�g����l$�l+|�� ߶�U�>n$X+Ѕ��g��a�U|��u�P��i�#Ybb�p�*ܠ�b(�����p�K?�6>���I6��	+F���~�YK�ДI�q$�����ř_(,��V�H-���5��$� L�
��yz�K�&�3�2����P}�����k����$ �!���b�m��Ci�x����0|g�
𶺄|�惇\uCj���M�?�n�Xol�������/p ҷ�:s�Δ�=�Xs�C�u���lvz�y�I�B?5��E��*�щ�/�	�6{Nލ�|�����0Kx��AZ��2V:�̂�����in��ƻ-dO"��Q6�[��lH˼K�BK�TĐ[#4����结O#�O� K��,���%F6t_j������c�G�:��������Z�\��`'��H��+>� ��X��^���1�-g�^�A���$_V&M9@���Ѡ�F����������x��:��ˉ(��A$��Cg�r�}`�F��ɧu���Mfn�l�"j�_����.�x�t�Z"6��n����Ҝc����D��ey�-�j�	9r���2�bYcb��Vk�򻺧����4-2��[�*Z��^;ۭv��@m2����,�S�DlU�M�[��lkI��e���}�OO]�x,����r����������F�pԀp�0-!(�3E:��1��[�c)Q��	��-�ľ4{y���e�v�8�xCFHz2�E#�?�jN�*;H8�K6_�e샮F�L���"US���p��-����I����Z�A�*��Q0��\"�*\+�ى7�3ց����2�S�Hqұ���z��P���[n��I=Nh&eźAfaԿ_�����6+�ΝǃL${|A�#+o�y��U�w�P��0u`�D[�Sش^�q�T9�b
����i��!Lb���5L�RZ/&����&��ӊ���x?�.9�)�0�5��*=g����	W��#�M\:ʌRu�KX��;s��.�2Sԍ�91>;&�;^,��Mc� �8*4�m���G`�ºߎ����W&��}2�����e>CK���O#bpp��QLm�:�w�[���f�<��B�7��kNtuF��	H�� ���*.���3��_��d;rXx�_~M��i�KmK�arҠ�Y���Ma>�*��2�>AO��a /���O����Pp@Y|nɱ��l���;���n��s�(��dp��Ċ��:p2�:ZxE2�����H��|��L���Z��<�`dO.��L�j4�g��<Q��҂)w�6��Ys��7	��ay�~؜I�C��@����C����rE��,x9��$0'Ee�K-��6��p�?��t�$�"��rus���� ��BnSGq�b��NP���l~��"Ӗ4����cԖ�A�0�����x�FR�q<�H�fx�c��MK�%�n��Fb����"̯��7� ����OE*��]��D���s9��/]�΀��or�
z-^���S�`q����J]t��]�;�KeW�^�|��\n~�8�%�j�Ś�	�Ɲ�Z�-|������=��H0X!���߶�P@<4��a�|���W���X��0��%�X����.��)���Uk�WP�v�_N{�"7�������S׾�F��5,jn��ZaT�к�6/�j�a�V|>ٿ#��95�`xj:t�B��Sa�e9׸�{�t�o�G&SN�)�
�(Y�^���)�h==\ृ�oH�"���Dvf�C�!���U[V��04��B�Y���Q�Xz���a-�N#�.���A�ѣI���Bfߡ'�XGE]�͡&�V�����H���L"8�$1Nv�����s�ր*4K@'Kp����mp`���-bhC��Vmgv��G^�O�;�R�9���m�V%�SQ�
���jΑ�2� �SI�����	ͺ��X�d��m�qD�{]��UݺL�&���%��7�PEHM���n��̒�.n���aD��ڭL/ ����o��q��8��Y �eb�JUl��ѿ���g(��6Q-��3��E�=�?8�L/��V#�t�`|m�I����7�u���#�ʩ괟f�m= a0<L��*f1���z
���4"ml��3���0��
ؓ݉V���^1#�oe�sv�������0Gt-����C6z �9\�O�Mo�������;c����n�xp�\���ݭ�s�_B_�K���Ԥ�HH_��e�p����1��u�x�F׹�\�rc�D�8.�=[�]�L^�ʎ:�������+o������ޑ����b`���r[Q�
��W�?�>n��fK��ة��-h�xW^�6j�ܓz��W����7���׍M���B�ˤ��"��<Jua5PJ�lS�����X��Z�\��X3ȣ� ����Zn��2R���X?�w�>ǘ�4i��:L�9=1,5�;�ct���!Qe��0x��
�)�z���AfK�ϕLχ�"������K-�A�0���ꖃ̸�3�bJ�!\Mj���P���zןYK�[�3�`�![/�,�F�8+���i��#L��L��h��%�f,������N�⥼r����9�����Z/�U�ʬ�[+J�`Ʉ��Wtw$3G[3�6��	B����\l��Y�k�G�W@ �Q��z�:,�oxG����L���+�/Ij1cd�Ƴ�Bf�Y柍H��P��VB�$���b���t�H@���s�ȸu�oa9$R�U3��t�	r�qW�l���c �6e���NKm��o�����N�fS����ɡ5 �t�%䢪9��R�"�F�O��q6���-��l�,�Bg��0�"�畫N���^�����Aʪ˘(%�d�n�-�6Ӵ.v�#��b���ɍ{��]���~e.R&�_+.m/@,8{�B�������`��W&�O�Ѡ������V���FU�.�<v�r'��p����*/�årj��Se���`FS6.��>��w��6��HH�ǢS���>��v<u@��#c���U<��=�\�wE[�w�F���1�O*'i_AL#*��A��;F*����*�}������2E��T�w�~�S��A��=qVA�d".ia풮3�!XД��g��,K��>٠� =o� �K�ބ�ɖ���k��4=����{ ��$TD0�t!=��m�����W������ʳ�c,v�Z�j�B����$��,�pV&�.Н�������s��7���n�`�;S�rx��ܹ�Tn�-�)z��<j����bq��pE�Mp��I�hJ�|��!T���I��i��N�X��='�����ئ��O��I��2�_�I7Ƕ��n�[�N����H�[tH1�5�!w�����ꠌȡ�Q-l���m�7�/ZA_�y���O6��������2Q�_��_�f���C��r䝕��R�:Ӈ�*��LQ���#z��/�̱�}2�C�E1�|�����D7E5Q�/˷�:��և[$Lq#������Gt�R9��c~"$R3P� ��hRs��O,%��WG>�~��r���p��e��.����H�P�F� ŎC��-	�1�K�"p��v�K#[HP �Qu�~/1��������t��!5p`M%��I�XfV���!�QpN�BJ�j
(��ɡ�.�x�2���	�t���jUy,:]�oBL���Mþb���J"{k{CS避�ɂy�M������uJat�WWIR�1D�Hg,�����}���7`l-+yE�.t����3�b><�E���ߪ�I�V-u��1������H(��"�M{5 G��x��8�G�37�� J��-���RȲ���!��НI���.�-����¹���,P�=�>��m��5���#\��@���O�cЛ�qQ�B��� ���W}�|BVQ羢Jd���	����ҧ>[��̗�[NH<�SBx�%��Un.�Hӷx��b��;�A��3[ >��r<+dWG��_��\����[�mN��_��ji�T�4u�:JO�ٕ�!.�����U^F�F�HY�K>!Gf2�zʂ��U�*�70\=���'�+�f��c�y����u��Yu�\�]k�,��r/�L�Y��ƚzON�y?_=����v�e�̛%��sQO!ܴ��鰰a!������ڽ�s�U��`�{�1�\�#RG�do�m�iv�>7y�a��\gOݔ_Zv�w�Q4�жM��,^�e�
j��������QqZ'�t��~S���/�F+�G��|�x�]�c� N]�diБ���
`�n��5ńeh���xVA?�K���8<p~���#�F ]ljx�kzk�9E��b���
��q6�ߣ���WV��P��M��P��ښ�)i���.���mq���3����wL~��('	�q�U}4��bٻګ��β��Z�q&�)j�
k�[��j*���ӆ,d[!��)���f�_T���4�H ���;��:fKC�jˠ�Ż'b�r��j0X� �KêrR����K*`��৐�1Ν�z��Y�)6K��c;����vE�ik%=����$��?���1\�fL�nK�~"|E�Tdq��q�ɞ�P��*�n�ɏ��l�.�(� ������5�� ��8��R�._|���`IvxЋ��ӱH��D [�E�]>/r����Ű�0J5J��	Z�@8(���V���ҁ�:C���;��B%�U8O� �tTx/Xm�^�ܝ�t��Z����E�%�l��j]�4r>�s��3A4��||�Z�o�_��h��#��{��m�ˢ�#_��d�����4��"�����{m3�-�3p����<���P ����/b��M-@ ��rB�w���������_w��؞����P�w��"I|/���ˇA�RV����f�#�t�pia��U�<ɥN#��'(�-E����1B���F��VUJ�Ktd5^�7d)6�cn����va���|M'g �)��v�%�t֔�.&�m�[cʒ{��4�#�֜��^,j���8~�H,�tdS�^
���CB��s��l�:=�&G��-��-و*�Ըdo^�~�Y^�E`�����f׋�`˲�\�EfG�kb���r �{�I3O|p�J܅��ԿR��RϖV�u�@f	�Ƿ ��0N�7=�!<�nf�k��X F�i���˞�4�z~�๐�͎��th3�}�%|�$�kh��6�Ú�2b�F���ȱ����
���1�{� �akԨ�+iRh�-���P��B=W]y��	q-���R�fR>^�mk�;�Ur3��y�_>��������A���Q�$�݄CQw�۬�ј�W,M��R�SZ�h'��A"1�qn޲az�
��,���2Q��<�O�kU-�'4�*�=�b3�5�N�Og�u ��/��#r��$�S]{S+�&7h���O��g=\���}�	�L���н�*g�uY�y����˼xv���Y�}�����G��lhӃ�)�_�B{� �@=먠��r!n��Ɂ�.u!/��q�f�m�p!۱�۱�+��y���a��ǅ}�4�١hs`<۲���\�C��i��$�DN��5�"��+	��E�����C@�݉�D\j���<y�_#4D ���/�|K��6A��~M��m�����1:���}�?�h��(
n\p�\gܻ[]�:�T�]�<�8[<`=!���!XL���=
�������e_A��#X����v�������D"�?�=]s���A#m�cn�y�VY��.�h]i4�w�JK b0��;�?[% �΋�����Ξ)~��g�3S�ir�A�����=@�,³���F(B�U.������w����O+ ,����M���g�4<��ⅈ�O�0J��euA-*]I���S�Ǭr:z�J)����y�Ы^|"/ԁ�7�l����dS����B�_��/�E8I'F�BaǗJHF��&v#+���|�<��Ô�E-ԩK1	n�ǝ_�}V���-V�cU9��M_B�['�I�~s���,����J��S�ꦢ	�>�U�b���+���wM��6��KS�om�OV�C��JƯ��~��![����(�y\4��|sU��e��$�BqR��A���輄F5tK)�fW��j�tjTВ��i� ������b���C����n�*B�L���Xp;�6����)����`�\���@a���tB����T2z7k��G������Γ�n��E�q�T����	�[�����i�9�7���2 *��(�\��U��S��*%���hhl)���B�S0����f~-�I���KFk�_Hd>���!xjtva�Ʋ�N1��HP?�7��l�=���D����̼�t�H,N�y���v�6N=��%���h�u����2U���'�m:�?<��R�;}��>��f�
��"t�J�I8]&��`�n[Cz�?Ō�P�쇓(�&�*aac�){IZ���u�L�ܪ������=CD��c�~X�&�X�q�;�Ga+�K�*�=⪊�0_4?�D̈ ��(���Gp�P��%�8'G7rz!��G��ڞ+![$NLR�fQbtQ"���®�#�'ē���}3�p=�Z� o����[�#MD��!J2�X?�O�cEǹ;�,ڍ�]Cm�6�2P����Yꊳ�o�����a����*K�"����tq>�o�{�gH@b��N� F}ּ��*��E��� ��ռ��8�)��ugQ�l�iYvW='.
�W%A�[I{��\S��mA�TJdQ
,���!��Z��Q,��IMR�(P���Ρ�K�*�{�������5����(�W�]b-�L���� U��m
��d�0&�;`e���+J��M)$`��j�N�"BQX�պ
�t3c��](ɭ\/"*��)�o��|v=G	˘�("X^W�w1PQ��i2�X����l�U�Q�@��I�������.W;�z�	�6f���ٿ1�<6�s��
?�sNiӳ��-,�\H�]�q��jp$���}s��([u]�nƣ�������Yp�h�*!�����H�)�80�i��{)m�*h+B4��^�Ԧ�*{#��Z�rU=�^%(��/ж6uk�w�T��X"(%�r��F�/؆Ba��mv��N�Nqh���b��<����hދ?���il��0��S�TF�X��Q�ϛ��ð���9�(�ř�1o���O,���BH^�����T�|�^b)2ۤ&�ٵ�!���3�}n�����~ܫ����T&O!�$�e��k��@7|���o������*��~ϞY�+��qMˑq�&�\_��?���y�;5NAˋ��ɬ��p�2� �e����jGy*v�»�&̢�.t�P��N�$�1J���h3�%�0���_��ۓ����9���qK��5�=>��*���4�T���(?}��:��e��xs<����I�+���r��EO%Q���2�7��v�X?����ΨP�y�n���Ts6`�@ ���Z+�������������>��3�	�����o��� � ;�Z�o]�]��%�Vi�;�o��p���f�w���$�S�7�Z��*f�d�(�R�x_52e�z?���'�l3��"�r#�닚�I

�^/��䂘�A�{?�u�zu=v"��rzU���_�N/UD��#�6���K���*F��FH��_�	��5�I�c��O��i߮:|�l�}��]��.�Yn(.�>�E1F�v�T��ra~~���7�ִ9Od7��X���)`�����=�8�n����o�b$h<F�o�M�-����;�@�mL��K-,�͉FY����s\�����+����Ȟyy�M��Ĥ�s�ƕ��:��~�h>��3�a����h̼�i|�y�J����kŦ��}]�ch�rEJ��a�ǀ_�?��L�TO"��zg ޺�Y/ ��K3H2����	�	*�qw��#(�hH�M�T�&Q���a��~-EZ\��Q��H��ʿ���L��8�k���%wW�l4�R�u�۳ׇ|�{��.l$�o��ȼ�/����/gU�hD�϶�l�I5�C-@$&_�']�܏�auj8��VA�TF�ۓQa�E�����[�6�p l�!�趿�mǬ��\k�#rB0J�ͿKIo�uX?O��w2�kT�S�Dy����F
}��zb��tRf�v��áF���en	��	<k�:������ψ�[s����+gA��զL黷��Qx��a�L2��*Ϸ��{a�̬S���֋+���߰�}z}���,�+E6�'�>*!w̽�Z`(eȏ��K Qˬ�~�M%��vPMZmH�9�2*L�T����Z,^����������r�Ѻ�3B68Ns��z\�j�IB�es�d��^�+d�ʡ�P���9YE���������e�&cK�v}X�y����8,O�Ү�%N�b�#�oxb���#����v�Y�6R��O���*3��c<צT�Z��! �l�ͪ_<2%�JJJo���'�{�v�brd�z���Kw�[Vg�&�!���� �,c��w�8y��,%G2�N�>5 !`Z�˚���~I������r��s}ᙲt�ȶp�v.�������z]��;���K�I}�n��cy�T�m�����S��w�g �rl�mu[�a���L�:�e��WvS6�����Z��E�1T�m	��^�|�+}�r"����7'����R��ڌG�����;�=z*U����䎆
"IV�w�o�?����+�<|Y{1?�GX��`�l7��Tv!���[2�U�O��B��F�Up�\��/��]�\D�ƶ:��1��t��Ň5]�3$���p��v��`�A�܀�NC���-�3��1i���Z6^})�,�3\f�ټ�����w�����%ٝĒ� t'k����]�eZ�<�fQ+=#�Z&~T����䒗YY��<.	��(z���.�Ք�I��;����y��`��g��1�����t5�#�����D^&�x�e�؍�%�E�[3]~����f�;o=���fπ9�>��z���� 6ĸIx5`̙�[���OX�I<B:'�=����Zs��ؕ��J�a��΋�؄�&���R�F��Q��RR��J��Ax^,���D�#��oF�ԁ[*�h^Zq�︒�}+-3#��<�M�
Q([h�!d� �������?7��/l�q���vB�Q��m�]���o��
��Q�;���RL��ɞs��֒=�Wr�S�5�B9r)]�l�vL<P�e�+u&��)a�Sp�&���#\��/��&��x�b��H����َ�xfaM��P�	�|�B�e-M�
�Zp2h������h�Dʹ�)c.�͏�mvw|�y�D�t�7�ћ��� =�k���A�43�����b֞��N\e�1U��������#�٪c���h9u�AR�R��I�CI;��x�Zg�R1}��W�_�@cO���s���X��nd���"�U���ˁ�kxс־��}���k#��d&['{ÜABj�� t_�@9�wⳛ��i�f���k���3̛-����(���fU����!$Uj�$YZD�D���C�ͥƱߞ�鑾��֒�j�W ۷h:^I!�H��9I��U.b!��=�!H��<����e+֯8q��b�DTu�ŕ�� @U̊�8R��x�X���OQo뚸|Q����Z��tF`ë����e-&4F�r(���(�8��WӫMJ�M��E��+n[be�]���o�Q|~qy7�[άՏ {��jK��|�
�ZU���Ԥ���V�/��ʼ��&\�b�F�[:�G<I{��Ea����	��'�R`C⫟��{�++�(��#]�*3hg���懽��ۤ^��w��)�R�y$%��L���KU�W�m$��S���onO��G\��)o�T��'FI���#@��j�>�����M&�K�63�����LU�,�|݋u"��ֆ*HA�if�e����=�QIB�n\9�_��� �~i��J�'�[t&����:Iwd�&j˪��v\6����vך�l=��6K��=!O���d[= fv^���S�Ժ�PuH�Պ�/�̪�S�!��~�,�G$x�\�@Ӽ���/�kށѼ���pҳb�����b���e�C���� ��W?��3��?j�����=�M�7Fnl��ݪ�� �o���`%����K��uʙe�z������(��H(MخH%R
C�ۊT��?���@J�y��淉)���������9Kw	+)�'^��>k���wPs��\��}o�V��RS6 ��bn����� �4�a�#з3[x��Kj�G�!��1l��*��Gn�������V�~�pk�BD��p��F���EZ���n)��7/���|�Nuz�c��x��n�q�k�g�Mg�� ��m��we�-*��A�熽�oP���R?�FQΘ�e���B��mSS��C��2/І�ۤAv�#ROf%ʒ���괴�+�̄\�^���L�JD�bK&y$ʐn�F�*C~m�wUՊ!��=2�;S��&֞�F�mi7�Ah�~7�-~3��xrϛ���ƍk۔.�~'�<
�#t,��K��Ymn����~?C�>۶�x pq|�ؐ[�͑�%�7�	\w#���J-8כZ|��G�{s�UwSxE��r8�ˮ���E�ܨ��%؜��s8jƻ�� sY��|�?ˋzW�����p%��Gy�'[�	�������]S�)kT���+9֋�7-Ŝ4�cB#�y�Q�n6�N_L���AR������O����ӕ�T��J>O���P��qۅB��|UO�t�6k�.͚�H瑒� Oh��W�u����m����T��D�r��] ���6��>XGz|>^��?CK1�j�M3����ȋh� �P�iJX�6窫�5����g�_Yߍt�dǬ�3$��%O�*}@�Ahl��>��%[��kjϑ�XZ&��l��I��E�
C\�&��>�x����S�G��]���pe8���j{%� �$�y�d�~l��1���Z�a-,�Y	`ю��{��R����'Y��Ѻ=��b��Iǵ���v5���L������"G'�c�3�dd�_u0������	9Bi��?�ȗ�{��k-���(BT�(��顢}��%�sy�VP��"��lv��r��ְlm>T���=�h��X�l��e~������4	x���,���ʛ���M����K֍�P
^�9H�F��nxë_=E�˘:�w0�_G��l�F���j��'e���g@���ǫi3P� l���stN��	�j<A� ��?{r:����ԟ��r
~@8[Q3`��j��˷?[0�+�wq����z���AL��7$=�|r��2M��֡S�tF����c܅�ggq�-��v����s�4hZ�g�@$z�~�+�'.�v�[Y�?����xQDس�P���3�%���u�� {x����m
MؘM���D�9�PD?�GLF�V�~��k��c�M��&�3��0�?�P�zq�����Ԣ�����3�����00�C:�1.fr��ӑ�fo�M8�_@�z���3�Qq��+ɔQ&n��yG<�������iqb�8���S)?h��N	�C����b�9-�voJ�T�k��-=6�X���{�E�~c^����H��=qz}q��ƻ�=�����l��깥1�ǒ�\�ވ��_8�aC4ϯJY���M̷��sS�An�ņ�$���D�����c44�l�Я��к,����(�i|���l�x�n�%z��\[��q��YI�n��|�s�gq}�;J�~��6OԪ��8��\�j{�mt�i���p�w
Qp�'�(���Z=5o��*�>�Ϥ�?��uy�  %�,"H�.:��g0���a O����raº�[�}9����ǣ����>���c��ِ�Z�'^"������KN+<���Q��85@=k?�H�>j+�4l5� ��Ų� g��ɿ��+�;�Qc}���V�Eڌ"����M8��5fm�)6�0�� %������nx(�# �P���q�d!{`k�.|q�*&0����	���yϏ�<\�߳�os,W�;��j�UrI�Z4;z��	C�e(w��l�O�B�@/��t����}5��.r���Vb�&�/X"���u��W��˲v����\�
�b(e9Eaj����hl�V�~2���k�'�X�wq�NGg�~//o�FZ���B�a���[a�$P]onl���*\�W��͕ʠVEWLgxS%�ɗ��,��z���T{K;fFįx�.����OM�s|)g��>�p2�m35��\�Y%�����S���yP~1W���E�1޸a�"8�EwʎҊP��o�T�h�����i��Ek���;����}p��*nJ��}Q�8�?;'=_�	�I�(nя�����K�`��&����l�gx�央R˞����Fl�&��r�Q�ܨҞ�ʿ��X-��m4���D33h�{uf�I��?���i5~�<���V?�.�<`g�L�we�"�E��*���a�"m���-����䒂�uG+�y�d��0�E*�.ĳ��<[R]W�mݳ:��Y�����W����TzWʌ��gD�G�
K[�v�.P���cnt�BP��P��V�,�M�������"��L6�a2(` �>y���p(\V��˂������*��N���N�q�ջ��Wƈ�盞iۥG�a<4,����%�a|�7�"�����k�Dp��d�=u�� ��*pF�䧕�@g�������l�Z��Y �
z��;���ɓ��sv!���e��t��y]�%�/T-l�� �ѸƸ>�9�ly�����ٹ�#�9����rԱM�{P���x��	t����H�P^7��W�oD�՘c�<G+ Cڪ���hC�E��b���8���+�d%�%'wD��Su[~�t���47���` 1�n��}��u��E�ƾNumr&�*��p��7��;>_Ao�D���Ͳ��z5S٬N0��@'�#�ʝ�C������x���Qd����Vȶ��?�u�79vwyG�}���mNk�	����S6��z^%�#b3�g��l-컨����Ph̑	��Aq� ������7�	4+��="�r�������oCI��H�`�_F-H��������i4����_N�*��V�U�V�_�(�>�Y�����/4�([�� jzC"+��ƶ��O?�����ˁ)�g0˕�" .�^�z$4Trf~��o�w��2*������e�1��Z�Z�'�b�s�d2��Wb���k00{�T�K�Ɗr!x��l��y;���a��L�C<��g�\�3�r�����p�?�<Q��f�;#0��F���m���tt`��)I]DrKv��0)���� �����T[l3�F�חC�g>o�8�h�6�4�oh��\J��e^E���S���g>�s&���𷠃�ǃ����~���g�&a_�ʘ�a���()WsAJ�v�;{����X6핲M_-[[��d(�5����(�������ϩ���yΒ���+�Q�3h:��>T<�Ҏ��/�e���O����h<g� 4�iI����a;Lݍ�p�LW�x>��|��v�	����"�[��UP"#��5L�8S�xs�5Z�E�J�̕�������(0v�����!#�:Ba�*�ϟ��7��������@D�O>m��w�����&β#�c_��o��v﮹:� ړ_O��k�X���x��)�m?�*G�����/0�5�~X��T�&M�"5�">��r������ʴ�9�iG`�h�=�� �*� |j%�~r:��x/�DA�=ּ2]�g8������1ɌS�I��)΢�����n���}���-�w���F���3�N�0��x���y��Q��0r�/w��^�����](�Nua.ep	�X���侃�r'��V�h�ćTIp$}���?U�h$J���{˧I�c$ϟ���&:ݲ���y�3���6��Sus�z�����9���ϰ-��:RR�K-'��<���F�}����)]r1tS���EZ�濘%�3�v�"a(^[Qx��I眶�^��TA�����.��f��N2��4�ꕱhg�uX���S�7���ǜ0�Qu1����B�K��m�|�s�a��p���Ē�����,��P�EI�}jD�5e���S4����t�igj\��ԙ��aF�t��#Zo��V$ �iV3F�J�]�������(��ss��j�G3��F*�����)̓��G��xx�����"�X�$��D��+{� r )1K��,jp����1z��I��(0��I���Ô�Wz��X9�<��9�ʴy��t$��}BԬ�L-t L���,�{��X(P(=��b��M�2�זJ������c�#��>�pgZE���睝W�.�-N7��1z{dP;�<뮆�Y�}唦�g�1��)nF�C��ٮz�dhx��a)�����j�Y�}=E��c�."ڀ���J��ik`��}Y����?�9ٓ���t�*��	�.�Z�Vj�Dl��,���q������g��x1�Ay�y��j��	,�B�_B~��4��h����v��SJ�M7F�Ǥ�V�mXqr����O:�hS�Ԕ8�y�	�6�o/�*��[�`3˧�&�������0��Á%���w�!!yb툈>�!�/B�X��?�?��[�����/�8�#� ���M�.�S	��j�;'���Zҫ� ����R����#�k�S�w��s�?�,�տ�-�{3�a��'��H�M�4�J����������u6qWm�tF��r�A[��~��/eq���o�=�V$E�gf��`d�(��&"�3ɿn7��3�5�Oc�E��o+H��깖��<$ "�jT�?�F�*���̱�}���;�<���(�`�����B�E#�~����A�XTκq_���<؊%�~æ%D>(%��/�+Ɵ˯�z�B��,^<��P
��%��%Хv�Xl��K��v_��D��bῪ�"z�'�w��Wh^W��|˟�d�Q�����3]�\��v(	C��B0���"����t�f;�Q�a;V�`zR$~�Y4w��vQ�:���*^>G>���Ӹ���Ay[7�+bw��B�=�Q��hT�'k`�3�'�u���#nkV��D�#������ha5�.��ou���Z���g��'>��I�Q$��X���x'�x��ԣ!co�W�i*;����$��i�	���S�M ��D�5H%os���ӵ�8g��8̠�����OIAp��Z���<U�B�r�yՐG=���@��
��z6rsq=Y�:�u�Q+./��Z�γ�␇{x"�t+�M�~7�x|�P�WG�5�����g��b �Z��S><���4��Y5R�����wP�w�i�;S!���m�E��Q+b�/B�m�f������r�����UD��9���/��Ј��q.ĥ���e
��W.�T�u�l�wm����C�*|��"zP�]����)@&�W���N�>�Z��Ֆ9F`v��K,b;���ɵ����y�bO
D�J�ʚñx�/�,��6���M�&���9�|�zA���&o3Nk�����b-�g��Kw�}�so7[��%��g�6�C���B�R�[�-�bc�K=E�ĕ��E>�b��|g�|q"�v�����؜���"��v4�+Tݠ���z���ŇR,�q�Υ㱞��B�+��d;0����j^���g_W�B��ȝ����O�	q�a�  ��t(���=I3�E�ġHJ�.����D5K���កa����B�\�J��g2Wz2��ލ{�*�3;$M�~���FvFQC���M�elo��?Z���c$���B"�hOj$�	�Iu�>A�wd�`�KZ/�L8�O�\O����_����P�P]�`:�s�P5B���2N
e��#~��T|kb�/gv�I��l����5�Vm�uf��}>c�0k�<���]�-��`�i[�S^Ō���(���k�`���d�M\��i�d�K�V+�����391��I6Q"ܺ��#��z��F�}z&����]�̰��5���}2�o���r�����וJN-y_�9�C�D�$63�����?�E�y��������X��X�m/O&��$1�o���ߗ��'��(Q�ߩ|�O�TD�0⸛yA,���m�ɵ��j�X� �r�������\oD�g�r�
_$�]i�+/ё�=��`��ޅ>A��D�șO{dz���{#�hЬ`�����$S(KO�e���B�\�y�z�F�߅>��hQ�k�Qc�����?��g?��8�!*q����IS<�>�N�B������wT�{'��~ձ��惷Qȟ���V'��< �6O���'R��[��R�M�њ�U�%2x��#�sy���,P�p��6�2����n��?���S�l@�TqʈY'/|M�����gr�u�B�t/!^�5���� {��)Mp��7x/��f����	d)�[�ϣ�oI`��}�k��NKXP�"����̺��O�<X�`qǨ4BZM{�n����j�]1S��Cb �0w��K+~[9/�鲬�p���Hd�d��X�E�K��J��h�#0[ze�Q0Tӷ��:'%3L�6�j�����-����S(��9�<����5�h̕���1����ߨO��/N?����&��#Ljd҅ # �{�C��ݕ~ա��
���@�/�'%N�;\���8�~�P��^��(��`����\�xx�vz�����O�&�В& g����`OD��P��O �n���%gH�x�@�]l�E�?Q���i��	d>K�r�v9���>�=f1	zbu1���*�C�E���ʰ����A��9xeM�sm���ƹ�#���@���u�?p�,�A��}�5'�>��ːL������*�PHZ}4*����Uɯ�$���ą���њ���G���
f�y?8���Ʊn�b�{��'hh8�C}o��-j=�l!}�?�3ld����H"
���m�k�w!�w��s��pu�a��������q����0V���hH����׊��vX��ʝ���J�0즊�9�5�WE���<�w�iO�Lr�ĵ�l��RO?��>[:�Z�r�;+�CO�4[��&���]�rb?d_󻬙�w`Y�t
,�Ywa9��!��z�(wo$����z������v/�`7���|���ru5˥)h e��7���<��Т������g��-��3�$�=""�V�Tǁ��5o�$�3ױ�]�pT

��h�;�Ua�-9$��#oB��ܛ�̸�T5���r�K��Z��uY���c��aH5}C��	����S���rԐ���Cr�?b��>�}���v��y�ʭ���n�����'��	��p�u��B�P����� /��-4�P��Ak�\�������C\�r*SH�MJ�b� � %[�PC~�oE��!g�~�Q�ࠏ?�����/���Ʉ�m�t��r
�h�-޽��f��c7�<��ތ�nm�Z J%�����L�*�h���`��xuԯ��uT.�w �z�|@Տ`v�5�ml=�ӄz���R��n�kE��J
��]�h�G�v|��z�>b��ݍ�	<�q�W��;�2\��^�!���Q�s�7�3�^�ع��Ӫ��x�qd{ts�)v�XJN�"���]~��d? �P��7��>,,.��S��s�nI0�atu��t�ЈP��)��p�V�6�З�iw[x��*� *�M��R ��Gk��|�
�#|.���{��C�oa%���鸓ƹ�Z	y��i�Xo֞�S��Z�*�2�`x9�Lt"��~���W3���d��9K��IWuQͮ�MIÇ>��}r�oR\�8��4<˒=֥ ���"M�O�u5�r�aa��J���0c�>�V��{J�VB;�Jfj�gSF�*B���������?^�������&$H�g�y4yH��,O�_�~�ܦ�Du�rn�=���mg<�/f�zB�j��C[$u������Q!p!�qc󭫙�(��8Ț�{��.~�L��nZ�;+k)}��X��iHN�S�ۥ@�+
�I���<C'���%�TnB&�T\�)ƚ��q�lē��V#�N<⫵�2��N���:i+��SsĿ��(���2:7�{���"p۸��˸����#�T9��Z�g�T���~ƥ�pUZ3x��Q1+¬� 9����D@bCe��K�Mr�g�j����N�B���ە+u�<B|e���(L�2�aM��
�@�N��в�iƷh1�ܟ.�{�����F>%�)�hB�@�1�����.˃�$AXC>����G:h�Ѥ�E��,O�:��E~ޣ��� ��\�3|�?�z'v3A�9u��ZԨ4?�}�����Mmq�*�@J�~~���t��A}h+���og�_���G%0SW"	�`O٦�d���V����=$�b���^HѸQ�r�<��n�{$V8��p:�;sVd�s�C/d�L:�հC��@��@;DkRS6�4`sIH�6A�)�a�V$5�C3r�1�L Ae�9�])&=�V0 �ˬ%y�T5ʽ����?�Z�2l�:��]����*�H9J	jղ�P���A����� Y���U�3J��^#~>��e����I�S�J�����}.qX9�B���d�%� j�A�A�$|%���vnw�x�|^�L�8��Dq��O]�U�b��mE�����wc˪V��Sh~ڸ��B@��O���g>H��H���1+��]� �fpz��;@6���2���0���1��o������k���0�a���<�/)�:�����%�F����+R�3��� {]�J�9��s}��a����~#����SŰ���Dn�T����K坜�-�%�v[2�t�EL�	�T��!xa�k��+��^ O/��B����Ŭ��ö7�"?�fHޒ�����׽��Y���.jvc�����7E�k�T�z9s%�i(���������v�9Y����}y&{s�Q�� o%*j�e+�4���Á��3�,FN�E�u�Jr�?!og�O�^�՘r<N���y�g����"��˜��8Y=�1]��6�4�xhk�SlR�0�N*ӾB>�|F�*���� �:b�6�J���
+�/�b}��P�Q�C ����� �N�ܒO�^)��6�z8�F�r�Ŧ���[`� X�a��/�p6��S@�t~���t�����>��j��KN���J;�U��
��Mu��R�[��8V-�����m�����z��cB������ :�}���Fu+�CJN����p��
c��Jܭ�7��+'�(rl�6��+�љ����J@Lz��]�6"F�;媛��(3Q=�����P�
�A����	
���x�On�ME�4���D��[ZH:7\+��r�t5]*޶R���
I2���aѕ#Y�g���Ψ�l62������I}Ś��Hv�
P�~�����"N�3g�my(T9�?�oY:.�fY��~��yq�=�H��)�$�8�	�q?���������:��w6�n�s�8H�ï��������I�|�c�������o��S�����Qd�BS��/�s�����5�b&�3�6#�U���A.S�`!Tݾ��Q�$ �	Nx����KtCb��C-b���6� ��W;n(�jU�;��_�I����H|k��T�:D���]\�d��
�fҵ�]�C=�Bl���&y���s���e�1�V���)��F`
Ow�B&���-4�R�v>9�r�^%��ړ�0����-�?g��6*������{8��P.eT*nAT&5�^�5�W��I�����|�ڧ�O8�(�(�0�1�� Q4��˖��E��ig��jRV��pq��p|�}0�leQ�o���=R�+��C�0 �͕�#e���_����4�;S����qބ��/�v*�)�>��yY�	�g�;��H��R ��MG���(^T�)��y�'�/A
� ��޿f�`��K��/���)�3��Cێvau��w�f�� %�2,�~�j��i=�=�"�a���JP��&wF��b���+g��_JA��^c�@��gWI��[�b��daY ���U�������!c��[D_�>���3���2���r�t�_�0D��`� ��?�^��F�*��/i���.�Vu����T��+ho�],�4�||���I���x��0�L !9ߙS}2˰9��)
�΀ܛ�塡�LFsݖU̎_�u�ߥD=��:F,����y��=/���0s-� ����do�i�)��|��|+׮����S1�Ũ��g7`�dy��`H���}p�8���{�{��=�~�#K���ބ�b�b��LY
851G��T
�Jt��}�6��2�5?2�A�A*�ʝ�8�56횽�U��.*�Ԓ*+�?�/����~�ɠdx��BD�������!9)�YHWl�����-EL�߅l��Pi|����(�p������{�V�	H�N��`x�#��r-|7�	��7k�#����;\��2�R0����3�ye��1PK��^���+D��3Fsix=:9�"v���u��0/��v��(��%��������ѝk#KuݐK[��ˆ��d��1�/�ԃT��Z1X6�|��Y+9��̵P;��.7(��`D��_��U}��2
�������b��
�f��'�JQ��b�A.�u�W��)�%ZH���';m��y� 1�q���_Cέ�-�_�x��p(�|Sye��"����7�h��5}<�iZ�����M�%��b��4*-{����-Y���1��/�̄m ���鍄�Ƀ<���ތEeI���a,p6�-��@����߱�1X~]ު!�I\�z�%2A���v]2G|@�����ͺ�̈�
�M��'�BL���1���3��a�)�ˍ�������'ؙ���ԕ��`����۹�T|'Z\�ӥ�~��˦��f9�w$H�M�uS�(w��*��ޭ���F�,Eiݨ7�עp9^}>`f��k����F>�����|̰f��bX�e���#�+y]VyȎ=0��w/�N�?��Gķe��`���HL��'8��zk�ZT޸I\I���h���&K�:�4~�YR�\s���ڪ�P:axDO��.�5��>Ho��d�$��v�B�B-|���0�'�E�ņW0����Sq��4���+u��Q�9O��*.�V�z��Β�=N6����s�`�c#6΃κ'�rhQ��֙r]�Sބ=(���F�=��I�G=�E��q7ִjΒ� ��ԽUBI>h<��y@,�ֿ����VBK��e�	p�F����<��z�g�C�WG� ��d�Ѣ���y?�U���]_�K����N0���#��=������= :�5��
W�� �;���/����1����j:��e�3)�ʙ�>��fq� i��S6��(d=�!2P���[˕�}JJx�i�o��଍��;���F�}�3�C��-P7������?��7{��T%�-��+�Bce���u��6}k��'=�gփ�=���s��_���W;o% =6-�D@�Kr��B����(#9�Wݢ&|1�\��pΘ�Y& 5Ŏ�ɛ�@Mm<_C�㲡�B1w��x�d/�	q''!�$��q}^���n�	k^�hP1ش�EJ'��.K߅�D�Lb<��l%8'����5�|Ir\7��_��JC�~ܴ�*�`գ�@�~Հ�=c��V��P�f!P+h�w�1������h��p7�Y��cͤ"ϭ+��?����07�0%i@�0�-s�ߛV�S<����n����1��UH�?��-e�6ܠ���3x@g}cmg�|�Tݟ�V�'��ႂ,7�����<�9���se�b�'@�Ʃ��л �AO�Nbk"��R�V�|(%4��NU!E���ʛ��!��\ ���$����d��bRVs���J)�&���EW��@���i���I�˝�����J*���l8�� ��c+�u��t��㢇oӥrƯ�.��ل���mGKE���'�O佴���א-xٽ �B1P9QXe9�fq¯�/ ��/�,��yeM x����(ΥꮺY�G�ŋ ���b�9�R�]#_L�\�!����!+ds��XB��U�։w��}�Oz_��Ɉ��u9��&����^��M1�S]����]q�{��]7ZX�`p�]L�X�D	Q5���Q���b��$V��."k�}�۪Q�>|yʧK5Huk���w����Ύ
�6�g�u�h0��%b\��Θ�G�� ���pɷ�id�Iԯ�����S��2��wPV��>M�E�|	rD.r��e����n<�z]��nN�G���K�)�O�	ۂ���o�|���g��hZ�x���:�F�����-�cL���'~�5�`��;�>�Z��;�,G0hM��~�^���l�]u�{���L̴��f�*	�t���}�O{�-g�㉸�L1����4�ݠv�/�»M3*��M��G��׵uz�s8��a���G*��Ł�&	z��'q�`x������~��	�`y��.	�J���m��Lz�D��ggPbN���P"��Қ��2k���ZNpb��a��J5B�>b�\w�c�}~ALt���p�gC���_��0m44N�Z���j� c+.��i�y!N�5���K��� ���!qMq{���*d*����&�I}��z_n�~�ߋ�||�S�/C��9�����=fx�d��l ��;���v�.���Ww�Y��,*�4�1�3��e�?w�N��r�Zd��d�����Q�Y�e���R�W �|bj�XAM4�n����\�5�@J�Y�cIЩ�{}��/<�й��!���g0�6'�W�U6e?3Xc�$�fX��j���hh���!{_g��<;� �j��N�A�Z�~�m��$oI��ڢ���U��mB'��.Z(����"b5_�L�93��?Vd��SlJ$�f0�m�n.6p+�/��>�
��_��s�{��n�.��Z��U��_?���2gҙ_)!>�Sg���`H�8{�2<2�u���b������򖄼�-���ي�Ŏ��Q�=Xa��e�c�%�jK��d�:���T�S���p6gdbE�ga=ԿK�q"��fM%~%��.�z��71�ٚ�#5O.�N�G������ay���A�R���|ӌ X�(ʹH)���wd���A2#����Q[�þu�qNp�K�)~�JFqn�Z`i�i�v>4W�!�C4�Q]�9�.{t-�|�oa�^��������Q?X����{���/P�mn`ü�1�9��ŕÌ���Ϩx��3�@�x��Ft�J������V��٨Cp� /�Hl��0���=��~1i\���WLh��|��<6�mM��B��{�>�f�U�z��0��?����a��n1�x��!��z6|X�UHz;��j��.f�'��q���˵��v��Qi��xS�eL��wy#5W9���A~fո.�7�d�%�J�����Z*�j �[ZY�ť�;��]R��1��>v�0Y|��q5NpGc"<��J��K,M����ƠM1"g���%�ҟX�ݓ�Mn��I|���*s$��X扳�����e�6��C4@fMsy�69س\K��g�4��c�nD�v��p��4ۙ��:����&�`N���i�[��M�,��Y[�q'������D+,P��z���'&�b��[�C\��{�V;�#+b�1.^��ǈ�D�^�ovz�{���S����s��|#C�6/.�W ��d�[h��$X �(.\�.H��Au�6�6nh5�؅Ϊ�Mk�	��>&��U��I�Q�L��vMZ�T��iTJq�ق�C���,�����j��](�d���Q?g`�;��g���gp�ɂ�'���-�L�q��1�Q�eL��8V�1��������]��0�#Q��B��'� H^oձR!�W�F�k��#�߻���X��:B�7.Nw7ľo���m���#b��E�C�h���!Y2S`dN��G0�q-H2�C×��r��ֿ]�9�|Ǩ�֬��/J��%@�_��NI�w��)�]n��><���"�j
����^"�W����t|�Y��/�e�h���gOuʉf(�ؤ<�H.�~X����#�?O)�g�k�����\�<E�05h�}}uv��Տ|��%R�{0fTHAC8�R/�=Ox��*Ǩ�1h�*|kft�ľy	`@b`���j���Ł��H�ć$�<{.z��(���2���Z]v!U�۴rd7�������˞�lt�]�$�_���s���3B��(����40ƯGԢ��N�>+KSr=8�*"��
�H�[T�<��W
���47��s/��e����ֆKn�
�4	[�F�N�&�8�7�[`��_mI����b���Dv���1���ta,��ʪ�;WmZF�̻�dziZ�
X�V�(;���P�GP�K�l���M�p�X ����ǎ�Й��gu����$t��tp�<ţ�C��b�!��h�ɒO�Z���=��*�oVHZB�5&�s��l�S� ���_�]J�=E%r���XDp�{gO�yoeQ��]ʮ��������˹��`~����ȕҵ;ٸ�_��i�d]�MJ�IY���#z]*�Ҫ� ���V{FA������6S�V��JL���jA��7��?�<�x�Ճ�����%��o=�I�Dޛ^��r�g!�"#�;)��4�E$셱X�A&�@ثe�g�<��Z�t/O+ǚ�c1UV�6Ξ����T�ylii��=l��p��p�BQ�#�1.�+�'_�w܅�Ȯ�y_2��ٚg]�t��yOH�̉����C���Ι?	�s~W�����IrKZ�H�ֳm��0�4q��g�Ƌ�z+/1�i�Rx�iB3R]�\������ߺ��A��?�rM�i���E��.��t,��x_�&�BQ�N%�L��Uu��g���G��;�&������#Z�u&��h2���=]�T�2
����=�9 �Aܩ�kM��n;�/�/�[����+�� g���̩e�Կ��b��w0�ZH���}��,�Du��Ͼqݎ�7�Κ�[�q[��F�̐Ǝ���8����M�ttu���#zs0����ou��>��i�	G��-���S%�+?I�������!QЅ�u��Y]6��Pt����[�6O1��2#��/��Y��틾���1 f��љ*���v������ޅ�{VA�g��
�`N�F�֐FR���~�wP��c憞��B��;�[���gY�U��ۅ^�ˮ8\z~ko^[ټ`��������js�����q��2�G͖��5�ՠ�r^e�Y�V_�[mK@�>���?�Q�Yo5�p �?��v1�Y�I�V���[F8%H��mԻvr�<nn����|�纫�R^\toۛn ��KJ�c�)_��b,�'t�2��A����~lʐ������[&��Zs3x}����OP�:�
S�Ļ�nA!�O:�9�]ϵf���w2)[%�g.��0�}���xP��@pE�{*Wg�*!w8��{d�%�e,d�S?6O:�뻣>$ҫ��kL?|�#9;J��3f)�ʀ�d㢮R�[��2�=��js��Eolu\)�+�Av�oyܪ�����p��-'DM�����y��v�=�P��'��EP��~��=�1~�K<��S4�Z��정�E!oQ�7:S�_�w��&����Z��re�h���C��Dj�	s�ғ�����Ĺ�7�{hN�sɢ�wŴ�\�C���I%���Mg�#��Vt�Z7�/8�|��ݍ�W.��&�r�N$�$y���`�B;�J��J�����?j��Γʞ\��K6&��>�Y�;�7Ц��E��mm���ѐ]�����-D&����Gv�5t�Nl��R�)���� x�����v�iJ�!*��Q�@B$$���4j$iM��V��Tӹ��Vi�*dm`��z�+�طVd���N'uK��V#�u0>��L�0��Π�H��!�@Ys�Ü-�<7�_=�Y����e��f�ۍQa�NM@��z���/�������ûf��Y;�4�3<�,rݳ�������a�ȡ|BYgy��mU��H;�.px�-������
|���PXp�r�d��^7��y������3���D��Eu���*�)���0�PE��B��֟���	�>����8�|����o��\�\����(��Rg�"L�� ������NS���:�҇������Rr�M�z�X4��]<�]۱��^8͉�{�tR�[-�3k��ɸ.��Ub.#�&Qrާ_ȊM�Fz}��z&�5+sa�E��U���4:�]�n�~��4���q�|�?U�Tw�c�4 ��6�n�7B�q�.�~��+�5G��Mn6���U{��!�T�luS�l{6:�Nm�tLi���5�k6�U;�~op�c2E�^bRP�U���{��H���ѱ���
a@2��+��<4�*ٍ�d���k�#�2��B�</�W��8Ȳ)S����w�k
+�ͪ&̌Qv��97�r,]b�����2���h��H!�e5�N"`�_	���y�`�>��<}8�C��ϡ����ˡ/4!v�}�4�C�٫�8��R�4�b����k��40#��B����hj���?Q2V��8RP�J^E!����3�;a{Q��ej=b���b�l��ʘ��)Ӹ��zݟ���z*���z��h	,�T�8��E	����_2��H+F��H*)�*��`Ҹ��\��m�����ք�����,^�R�B;������g}z·0��@([7�@���(5��?�O�{Ym��~eC~�j�m*��t
U����P���F�Z�#,��O��� �ea���ذ.$�r���1q�S�<H�.�>d������Au�H��ysaأD�kR��x3O����q8���y����تZE_����0��H�
��7:����X�X��f�LIj��u���*X��T�$[/�7a�O0s�t��L����VW��4�ua����!.Z2�9vX�u�j���J��w*���EȘ���g�i�H�ra*�}��ca!��z�*!b���u��4�|l�oe���6)�O�}K��;En�n�P�/�18l�#]�_�\l��R�Uх����}�`�\����W�y�
�T�T˂�iY��5d�s�,�.�7�Hd$%�ԃ�QN���'I��X�e���9Ô@Qa��W�(�ޱ�L]�.�B��%���%C�G'��-�z���zVc��nDC��`|��
d��R�r8������|'���ںy�k+fWW6�*�� 'i�g3 �!�< o� �Բo����~X��dVn�J�pg��BX�F����ߋ�{�5��g��Tf���m��Qٗ�,�ԗ�dbv��l<������ibZ�y�"<�4�{�d���z�R@
�I��!{�Z��*W��
Y~����Ji4���{#�z��&� A�J�h�>��R8��4����a������'e:*Kx�"�2ߨ�zi�.{I�����\#�W�+wFO W���{����!�KQ�	�Gn�pCP�O�N�I��$�Ch�R�Ǐ����S����?&%�'�<� �N*O�����詳(m�����l���̿ \|E1O�ԭ��t��GCV����>�	 ����=tsC����I�q/��A6��Y���=ro������'����xp��uSN�^���wЁo=ؕ֋�ȿۉ�*N������AtyG�wZ� ����d�CY��ʩ�^��^���~O�`�<�Uu|IH�����z+q��p��GpH��,��o��)����jr.�{�� x��h@�ٍj��p("�,�::�@��5�!��ts��g���b%F���,¯��C�H�+R�Q���у�m���wd(�({V�|Y2���[�wM	`��G�`|�SE�`(=	>�L�������!�|c�j�.��.�j��b����K�Ɂ��M(��k(���jB�bZf���K��f�_@%&2X�Z�#��3�H�w�H�߬�>��|T%�����O��,oI��;�nl��
*��V��)}{:��="�/#�"쩔bn��C�v��>u��:<W� �d��j�G4��ǡ4�O��͙�`�<�bs��uD��?�yJ�t���m5��	ݜd�]m|u�͒eh�'T,i���m,.�]
����Jq9�O��
]�I�����e�19��`M� V�5vd��+��E���B�2�@`�x�i��S p�K�Og�E=e�-|�'��E��y�]�9�R-װ�D�HZ��^cʿu��e	��uwS�H8޿#��y�s_�ڝ��:q*�����(_�b)�P! �k?�r�k��Ֆ|հ��Sᢎ�^�n%w�h�P�@�]��ލ�q&�Y��&�Ҋ����'"�s-؟���(po��+��.I�A�̸��P<��8�4깱����!E�0թ�j���l}|���Á)�-��/kR�������c|�%������ Z�flD��h��^�[Z��7?n�l`��Es�04��̑�L������|K�0�a`��f�D�ߕ�< ?7F�� )��D(ݪJ���N�>55T�u���<��x	�q��KS��c��'��Gv�t|(v��ۃ�$LHG�"�@`����˦�Ͱ�͐1u�M��ʌ�*��ZW�a֦���r���ά��J��
�.<���贝����.N�a�r�N����8��!���1��b,�X�f�m�,+v`wA��2�B��pMiؤ���)�*WYRBrH?
��x|s��8t�~M���E���U�'�X����V��Sz;`ׯ�h�_
������?j[x�Yɫ��A���J7�<,i���-�O%�g��)�81ͅ��n_]F��c�� <�"�27y���{�)^>/��I��:+�������ʻ�y�ʪR��	^�Q������=�cxJR8�ȏ3\����J3��6�';K�����S]���%4�c��11��H��p���@��r�:�6>�4�/R���_�zz��@_J�< ��9�hF�������N����zzpk4+�"�kf5�Kq��5�>��c&�,�^7�d���/m�o�:~�^V�:T�j2C�xo<�{�E��Jb@Ib�+_���[Dá�~��U[���2p���2D�-!��50�ϕ�V�^���5t`���ɡە��OY-*��Z��0*�G	-�F8N���m��a�ڈ+Z"�����\��� �~�(�sW\3�}>���XD�#z���=���3e��O�7���^x��DE��U����P��!V�dI0����`_s��,-��00o�������M���Rs�*�w���U+H���*��
R��{T�sTyO�㌷;g��NF�=t�֗Xc����f�Ҽȟ�.�PJ����Pc�w���)�w���e�5�t�?p�ZϠl	{d&��
B�O�����)D��W �a]g��i��^/���d6M��wA֛p�I݁q��%o����t6s�h�̘eT�}"e��&~�nz�L�h��M�;iٛ��BO!�Bf��@;{\����2cw�T���Z%_�̸�ˆt���e�p1��{+qH�z�%�sX�j"��bŏ���ؔ��6�P�+D峦���5d1�]ˤ��6cS��P���l�Ǭ֢��.�${���w5V$�	K�6����[��4KH~�?��n��zA�2���\�/������.�K׍�l՟��:A��|�����9K>�0ά~,I��gqg<�#�a����)�4�ç��d�C����K��)���"bx)�'p
�	�#<�rX�_�^��$�1�moNi�
�p`�Pt�SV,c:��}�'r���y} Jni�΍*ꜰ �Qr�y�)�����{U�ҫUyWi���[0�Q�w�(��x��f�!mW�����((���'�T�!3Q��Om���`�{5+{tg�_��}8��I�
�+`������E�}*�k��z o[���=7j�d�/3�����%~�P����\��EU�d�h�n=�˵a�4S�lݦ���n�y�N-Z�P ���)Ϊ��T���y�t���-��tjw�4�#�kԩ�u;ⴾ,
~yH [`�ՖLM�r���o�N+����X"���;y���(�&�1rp0�Y���0��c�%V�lp�4Иl6� �9n�gi�돓��1���=]���G/�>~�@
�����"1,��b\�>5�^H�j|�H�^�Q���C���'�p �SR�X�
�%I0Cwlҹ��[��F1���k�ky��9�,,V�Df�u�W :�R��haD}��
��%GQ��`�(͆���}���n8�p���P���	��g��v�q:��-�{� �,VO��?Q�j����r��oe��s%��^�"H�����O+uN�)6���ߪ[��G��UYۄ�T�sn�
*FF	��zY�����E@�<.��=}��8��_'��}~a���G�R ���=~�@#k�*�Θ3;��s���a���9)ig_��6�6+BP�`�	'Zf{�7���'�9���t��wޯ�R�|����r�K+J�b��T컸~�'`�mX�Wı�r��<Q���ӣyUs5��-ɷV#~3����1����W	��o��Û�!z�R0���ː��b���_��A�hzR���ׇ���|�q�Ȯ:���	8E�RWi)"	��z��<�d�T�C��<S�kf��+�%�n2����\���u<1ɸ�Q�R��#�ȋ�_nu�D�i��V���í���/�|sY��D)H��v�{�'~��
��jSIf,lc�!�:l�9�FB8�z4�`�@��I�u���l�	����8�:�pƬ����^�B�`{TbX���s��*zwӚ�WG�0 �𻵲{G	���
���tu	 ;�2�j���^7՝*<�ֻ��ME�F
�e�1�V�.�vd^T뺈�ǀH��l�v9|�ǾmU.{������'k�=��L ���r?U�����ݮ(j4��ޙd�A�lĒ����)�rT#χ�Q��)���VZ�LѼ&�U�/���	oRE�Ƴ����0�B��Jԗ�$Dot�<HxU�ćOuѿ��捻M�X�G�dU�8�w���Z�8VyfYk�k���j~�g��݌�@��u� ��ߌ��"���򙏶?j1(�Bm�$��z.�1���x��؎�Z=XM��S:	y�K��l��zM��%��]��\��F���8��S�(
��'��Xs�/o:�^� ��c��hr�h�sЊ�(�vu���?��茔�j�ɯ��ޢ��7��FZ&6���fVD��N�zЂve{����˗C��r�i,�`>�Bvy���o�=�%�G �6��kT����L��B��\V���:��+	�6[ ��5�Z�F���k���'J*���y��ǳ��+<Վ�g�aM���c3sfE68���,s`!	�
mC�8~������z�p�������m�����y�d�P�v3�c�W�^��iR�'�����=��F/@�D���^sw�Px��(��R��Z���cu�L�xxؼz�Cե��!�;Ð�������*Dɗ�/ꨠ��{a P`�����ؾ����qͧ;�c��:]C��U/�b��x������5�vP� �!\0�h��)9.�R�՜�meOTS���r��`pQZ��"7S��\�<y'jGG��c��74�
�j6�n�^�-)��
�TF�����Y*�d��Jqע��h�_N�!�Uې��0u�'ӂ�x���-�pb���?�v[�x$FYꘆ�=$�LȎ� D�b�;�'�K�[g �e�3�<���wK�͘ܛ������L0���0џ���_w���j�)�O�v�Ys�?r�|�� Z?y�פ�����D��%�f,i��|��-�a�M�W�}h=��f���x+��Td�0 ���-l�E�ke&=��+��Q���^�I��,s~T.K�qt�]m���Ҧ��L�QN���/z�	���jZ~�k褄����u����Ve��H�%><6��<	����
HA.5ME>*�t��L�+͛HI���:C¾9ͬ2R�v��j3ؒU� �qA{t��n�=����x�q 	��9�
�6�� 怳WҖ-���w%�"��xgl-3!%(zo�>2%��:�^22 ��h�n��^\�e�ժ{>[��W�w�u�a�}9#���3�1+�ܥ"�-#|Wݚ�.�2Q�]z�۾���i*O��c���F��s[�&q*�t
1%�aoA�R�g��d��EG����YH3���7z"�����[j½�+(	O{6�e#�ʑ���ñNﮝc�=�EL�xo���=��	�����@�޲OU:&q[f�"����c���y���))�*!�&?���`z�*5yT���	Q�6�M$W�N�� �o��4d�W���+$��ŀu4$�8�^nm�?k얶���|��xEqN)tq���.�՘?He3��a�Z��"m	�=/G�� ��ƃ��ޏ�X1�B�x��=�z�������g��d�,*��!3e>6I�U�*F�ߓ��;�O�����|�Z�+�f�C!/��(�g��#�1�|��/;����ڶ�x-�"�,�f��mh&GwpD��9�!�kT�ޒj+�U波[�r�݃̀�B�k��q�S�[���r��\�[^�`�c�g��!����
���pg����2���m��g㇋�i��k�D��Srl
a�O�ˉ\�M���}~��F��{�\Hxp��3�>$�j��-��y�ʎpƽi:8W�PD�p��X��qlt������m�#��I93�\��Z���&uꓗ��I�jm�*lYS~F1t!���ic�p�R?�� ���N�`�B���,�<���^�RB�Z�fS��� �-en�:�8�Ikk�1J#}/��D��^7���=va�+�9:�:�,��i��r]w6e��OL�]��f���w� �*�	]�-���_Ǯ�����=Mvc�*�&��B�p�C}��+e��|��Wlt�Q>]#�J�0��3���Q �qm���bhg�ꧣ�c�oˇM�r�-��\L��	vc�M�Nd��;\y���엖�c0+�EܹB#i��$3�=�f��7؅l�ˈ�� ����}',���c�`��&���3�P։�4d��p{z�'��!A5r���#pq�J�8a��eNT�m�e5G��u��I���K�Y-�t؉ 8���C?]F����Ϸ*�
��q*��hC�#$�A'�?h�Ti�P�'Db��_DVE������\$�8f����Z��o�{�\��\������]�_Qϲv�!yi�Ee~�H�<�Ou�/e�LS��|���Ȝ-��R�<ޙ����5:�k�W��).b$�T�||�`��H�3��<��p�
3����<�.p3m����K��ڔ�a�	�i��l�K��2W�VC�!����wBbI�Y 9�������o;��k�#�l��U'���E��z�o�/�'A��V�	��R�vz)���Y�[j�kNu~�n�T@���%k.Y(�v>���!x8��F5EMT��h	_]&%d���ϗE�����/�M�m⻧��ش�]�Af��K�� Gp���@V�D{�w�~�י|
E��7.�#�.&Q�^!Q᪠���v����^���Ի�����K���>�?�w��hY��U?��7g6	�@ٳ؋$�c[�V�Բi`��:~�i31���x��Qsh{��s�q���mL�;�9ܣ�n�X��ȩ���cPkC��C4���R��g[��c1��Xƍ�	$��1s�>�p~�!�ԠU�u�O �gj9���&Fh5!SR6��za�s �4�(�B�_�8=����Y_乫s6ES�����݊�b6G�H�� �C'��)��u�23��w�|�oa�+V���>��m�r��%�U��>�B��m��FI��H�4z�1XM����w���K�����m" ���cO�r��]]�W���s����P=�!C)�Q�G��<b������*� ;�IY�X�
l��n��v�a�=�2��<��o�zȑ7��Cm��gƿ_>�|�HcX�ޝjV�ZM�a�Vo���%�g���-;W�q�|q���3��3��2�.u둚��$><Ҕ�&7g�H,.g�"ڬ1�b�5�P+
��<��Y�He���V��!ǖ	�8QmA����UH���_���I�R%l���q홂�~e�?���ޞ�E$�D��aYmd���]*��?�Y�|�R�_�2�mNr#$(ͩn:�t�ؕ؎�(){I���B:�3��ѕo�m�m��J�5p'��~�^$p@�BME�R�☧���{���}#�EE�f�� �sT``!h��'H\���N-u����$���s�L�ާ>u5������k��kN4܀+��1ܣꃫ�=��#"G@0W+��m��U~���Le�o'��0ˈN�G[X<X�ɐWdt⭗'2�*jx�9�g"����1H��*��dkޗ�l��XK��#΂�!�W���U��ۼ��|�ڙ��+���<N�4b�}��k�o܋����� �0]_6���KZ��[��4�f� �;M�����-:�H���኉�Lij�93ϩ�3��yA
����i����A�d@�z�-��*@�kx�{��J:��1�w��ţ���d��R�v��5������Y�I�)��Q���я�z�yW�d�zPN�|��E����&x.�H`f��7�3D�S��y��J� ��"ؤ|�E�)�o�	_<���f~�h.��g�y<2b\�3-	�w0�S�=�
��O-��ڋ`P߾j� �F�MЁ:%8��w+|8z����b��AT�����'_%�Gθ^ c��&���ў���;���l�'�h�=�r�e��&ߋ���6�%��R�Z{2��'{��%�C�Y�jT���T�Fx�t8�����S�H��M��!��6��j� Q:�ONv,0���u[��~�gR���+��b*��2\����P��^�ZA$�s�[�|�x;��^�ێ�u���2r�gr�\�L|�:)�j`No��R�2��y	�󧻟���$|�аmU�{�S-V')��zL�?�N�%�ݱ"_)�	��p� �1��f,y�scSu����Sy�G��Ps';d���<���Y��1,g"�I��.S.���9fE��p��Um�8t]84�ɹΕ�F�Q����D٣B%����L
.g�S8�A�"���L��"�u��t���ɞ�9� ɺ�h�A�+�sClՋ�.���(�(q��I��������/�K��
~Q�%|�2�C��z�S�Z;��c�EϤw��Ͼ�I���#�%KT��_/Pj�,zW��?�l�?i�Q͂��_�c[e�v ;-(ީP��){)8���r�L��aĤyK{[;�[F�X���RR�SV���}��*p�F	}{ �%lX�N�?�ǜ�u^�}]�#T����پ�2ؕ��q�@J�2��ug��,�4J*c��@�:ˣ,�\Z%;�r���V8�'w����VS�C�y̻��dKmZh���整��Yi�?�6��
6�7���=�,go�g�x�?|�����AMVjj�y��/|�-V�2�t�Hr�r���j�9;��q�#&���[}�o6��ec��عO�:L _�ۤ�5h8����m/uJ��BB�L S����<�%�֏.B�k~�ҙ�6$ͬ�P�"��>LQ㜼���'x����h��eY�����@Ш�e�U��w!��jujW�wa���J��	is��r��-�=���TE\�a'��0�y�+�=a�4*�.۽w$���M�<��N�w��b"� {Y�^�|��u�+U"������ya��
 ���u�
5���=����#y��/�?��}��l E�f�g�♌]�dQ���op�q�Uz=������yxׁ.Y��6yz'FT嵭�]8Va�>`>/Z 9Ğy8'4�G�e-���������XA������j��oh��+7���Bˀ@�X��3kfƇw���Gm�3�4J$���nc�?*����':���O9�B�Bڊ��Y5�d��xM������ڿ+�\u��I�5��}�E_��JYa5��SA�g��� �+�+�zp5p
�\�M|m8�����c��.��ZV��n��.P*\>"qp�9��
�>F?)wY��u���i	�K�)�z�i2Ccw��(�Nfv��T2�}|�:q;HT�2�8�H��"e�M���,�>�A���'Mx��CZ��!*�֏RSv����7�=9i�-�yՠA �
�6��rI�d������*���`������j�8��.�]���{�mh���V�]��$MxZ��]���u�K��p���p��*���� Zq�C�cHO�3q)��H����qt#,W�1�� 7a���1��ߺ&Q�s��)Y��W~舐�Ajp�q��6iȄ�q�N�xpq�ow�o��;�B�����G�:]��GL tŴ�a�~`�(7(�'�'�q�A'���0�\�Y����֒T�����oܜ_]��eJc=m�'#44uP:��Pa�2囂�
 !���b��+��>� i����f4s�F�*�XYP��Hn��t���q�hy-�J�`��2GT��)+��_oAM4,�Xu�f=K:ʞ�J$X��_t�yz}����$d�D�*��������y�P�3�3����`�����7�P�o#�ھ��	;�	��1���^�ޖ"O,'d%�^��i��i%�+%vZ�e��'+qAX��4j���Rk7�G�3f2�rK�J�)��aRʯ�EZo�������u�VP�����	t��FeG��<<N)�	[ߜ��	TPZW�����C�h�_h��}7�{s���C	�ܨ�-�1��rCX��x'~����5�ra�8�옎SC'�@�����a���Jk���;HE��v%�	�0+��>�p��FJfC^F+�2�#�v�������_���s��1"v��%�mB��-�V]f�l4O-B��ٟs�R�O7R~�.I]��d�"�Zr�����n������!f�.5����e�2��	�tLD���懖� �򳅶�[xE<9`��)��xg�	�4{AS�
��2�JM��[Li\@�a���&�T+�|^��Q%�숸w���Eؒ!�Nm2�T�QI@�ʘ�c&��(���F���;1�_c��
�ΰ�i��LCTy��|���]���N�ͧP�$���!��
��v
4�(��P~���{A�	_�W#O�d����_rS*W������|��\�+T*j��L�.�~�*���5؁a�Q����X3���I���kH�w��3_�f@�}����i��-�� 2��ڬ��('.'��?�����f�@�����	*��g|�@M�!�,��j�ZRos��m��O�v�ŷ�v��z�����ER`��e8���R�8��>��옺!vsݪ���;��&z���6�4�����F�.��!��Ua�߂��@��m���;�5�r&�,(�$rE,Ny}t5�K�`����C^fNܚ�4�������u�e�y/!=�S:A�z(�(Ĺ01���]Wm\�̕����V���帮7(Y8����2����o�*~3K��4��������S�'�L5(��s_S�-�:l�r~YUS�xr&wT(�������g��Ҁ��R�s���}���[�4����V�㆑�䟺�� }W�8f���Ǌ޽f�2��G�8�����'�Ɵ�KXW�C��ҫ',���d*����]��'�!��}�Ė-�`v��by;�G��oq}.��/!���+�$}~��n� &���~��
���N1���G&�ϳ���c-Y�ȑ���2��G��ʖSkv�`�#��UA�vd�,((X}e��8��N���3?B�D&��$�Y}2���QHhK�g��i��r�PƂ��
��K|7 �p)�uy|�f���7���יc�ش���r�F����jJ'�8�Q���PM��\|�P��a�	�Ң~�|��
A��dZp*��r�d�ܣM�u&- �`��v�錞ؘi~�7�Pr[~O|`l�~Oj'
\Li{�7�ή���mgplըsT8���-���O��+�GϤ"ČQL0��AG^�M�l����D��P`be_��fm|�~<����@`/ơk-����Or<�|���*=j!�+	S��%.�x��/S	�G�?�� U�pJ�a�ri���6��6X K�
;8�����t�6���TR~��Z�m֟�;��æ
�2�I����]���[�P	��hӨ���f�S���+;7���X��:\I��,j6~`A0s��	mX�-��r���8m��~���5�Ӷ&�������M�ZÅ.k�y�>f�1�
�hp.�	H9�1��P��C�o�߮4��3�j`�����]�����m�vV��
����%p|�Ir-w�Z�nG��aN�ʑkh�}�|K�q
����0�x���Ձ�ϑ�*�7��dN8	NP�*�o�)���C]@R*�Bn�v�#t��_@TqL������������/���:�隈�X%�m0���<#�=zg[r7#�!ݫ�a	cv��������K���J�yM����=����I�XF2U��}�����W��9]�.}.pŉ}�O��(�����.�^�\� j��V�k�lm�=J�܃��N�Z�Kb��/Oz�����t^C��D��gkD�ݶ �?�d}�|�#�)�u~��DNp���kmb}�/�UP)�",2��-RYD��J�c�k��!B�D&�h�a���Ed����A�u
�>�f��(��5(�K���3W���Y�z(�dG��X�3�|���-K%I�1������i.V����4U�b���"���5�O��ݘ/��yK���f�7ܐ�#�/Z�_��#v�]��\��mc��wB>P�t���5xQ�v�B���Րs�zLT��]���
_���,�Ś��2��+�c[ W���[�I������@0�F���QVVN�ŢF�'b�^٘i�Т�[RsI��|�%��kS\?#nE1�˝��;^�?���Q����0�K�-�.���YDCۧ���շ]섰����b�e�'�̣j&oğ����h�V�a9� Ag���>���&B�L��Ir��f����B�:�#i�_�?!3d�������v�.�W����i�3�J�����A�(�_�s�E���rQ����A�s+N��ݴ�&�X6L*����y�}�X��#%��2􃋱�M�m�M�/��SpM�j�*q]7,�����q$�i���������IZ�Iۘ�V8k��;#Y$w�O��C?��3�:̗ȓw��,����E2��35>�k�p����,.����a7Xs�Mg3���� 0,nAM���e,�8��t�>��� /�B�� 峰�=t���h{n]�~�5�G��n�F;�q�������Ϲ��'�D�I,Nw����-���;���� �P�����p/��������N�U5�QgT���X"6��k�1�4l�JSOB� c�_�1��e\�c�ID�#`���� ����xF��R�b�__x!o�����} ����3M�u۰�`WG�B�;F9q�7�3������l��I��
{`qo�Ӿ
�9��2]�9��l�=?H�T�	�?B��,jX�Mw�a"g����A��QL\�ؔ�p�<g�e�2�E��3r��	�z�v�KE�/m"���~QB[0]�<���t�&M�hvDp��:r������ꅌ`t>RFz��z
�'\�^��s�!o�8�8,x�ETq���,נW?�-,�T�&��J����H�ZҰi�K���� ��{�5ߕJ#'��������^����;���v��.���G��8YR`�b���!u�6-K���e4*.�(�%:���hV~�0)V�l����PoMut��\/�@��A)g����{��!��<͏26;u�}����;��!͑"�C�.4Dgi:h�7�/�W��Nw��#�O|ݗG�<�w80�}�gc,A��M�y��*~0��L�������, �F���p]+G��S��݋;ފ<��~�t��8ߌN��j��M��hWT�> ��`J�nKH\�T`&�,�����d|� �������3�A;�L	y�FTNH�4��5j�8���[ӈ��~��Z�rIV�6o�S�,�ƪa���ً���)V���4�F��J,�?��Ti/�t�u�G�NR=~��t#q�
���ơ��q�QKϧ	.�'�~]��LQ%'��m'��]�>��Ґ~������Ψ�Dz�n_.̳����23��vv��B�a�4?H/G&�GCm�κ�/�kH���2$�3H�V������C��7�.G誽x����kN��ɇ�)����ݐ�,s����}b�[�.f�5�-��v��zM�۳�$ÿ����<u!�x�NH�޲�\��1��a����BDm�5l��"�K��Ej8D���0�/�tJt٥^ T�)`#r��)�Lqm���Vx�V��,-���ur�`�Ҳ��御��xc]��[���ܝ ���W����-�2{����"	��R6�7{�!��T�]�W%ԗ�D�9VOY�o�c
�{�Z8�bd����w��T[��w��ŷ	����jP�u�@-L{v��K_AC�P�������ؚ�z��W}���� ��������H�Ĕ�T#lFMXԉ�p50w�_9�/U%o�K�1X����N���_�]Ӡ�J� a�0H>M����SC��7��[���P�,�bjR����]<���n	����7%���;�^�O
<��+�r��F>�����&Bt�Y�	����	��ʷ�*�f�1'.#�c��Ƨ]t�M8=K������n�w)#����k�N��Fa��k�t�y��Q[��XiPc �G���$��p��v%�^O�9S��-� �+������.���t�R5��6�&&[4�T��6���	㔙�E�t����t�{�t6��W��k�ȏ�_�G.7�
��&-��>6F������J�����N�h�~���ߪ���/՜ۛ�zk��o���}Dr�%���|�T���C%)*DH�B�%1-D� ��v���J�I���"����i��6�^M�L�̃���Hb��䃔�ef��j-A�YC�B�֘�ʻ���g���z�N���q�-��L��"ZX��Ϸ��DIɄ� ě��X��"x#v��ВpR�'���u:�n�W�ٰ-I�:�V/�R�ܜʸ�Q�z~"�>��6�?�8�`��p���1�����ȍ�.��J��z�����OCeM-Ё�i��3�/���2i!��r��������?}��`l���M�w������.w�0��m���_�ywP�2�h�7�f�#��|�2\a�{~`��޾qR���_F1[̉/} ����YQ](Z�m2xl�Ae䭮I��L:��ݧ�(U��J����������H0��M��y���_�^����Gw����g8	�?j��oQ�����u}�?h�٭���:�k0iO�d��^s��^�� qU�Q���'P'@�^�� ����x��|&�8L�)|����	*v8�kg�o�.���C<1���%VT-K����*��iv��?��yY��v��S�G�K�?c,ǡ�2��6
�{Vge�K�Տ����z�C���(�/��R��x�l$K�Ԭ�$�@�3ۅЇ"��Y��EՏ��V$��8r�	��4��;�3�z-c'���Q|�w/�bor)֗(#qɧ�����-a:�����t��ֲ���]����v*s�<)����5J�uYy+�3���7�>�]]j$� m�i�"���rm�ZKmR��r���z� �X-A$��R��$�e�*7/J���n�.r�t'�o5\ܪ~���f }w�gU������`-�U�}�j�s{|�E��v��D8�{��j�/}<�N~)�l���dR�>3N؄SN���O�p������ka���I�|H���C����_
^����qHg+��2�[@\�ꪩ��܎Yb8~^�i�����?$W�[(w��ig�l����7�'�\`��po�`�mɋ�f���2�XL�� �%�P
��41A��v��)e?���?���\x��c�19s������]�fVk�`H������b9���8�N��y��M���lB7��"9A�b�/����iY�b�ρ������@�_a��@����P�VbyVf'�]6 Vg�������w�����C���G͇�)e'$�HB�ͳ�n[������}�_���U��O#q�u����R<cFCY!�xO�1t ���c��"���Qq����֭���
O�+��ט��Un�$�MG�����;�J��8e0��%Qe��C;D���� V�MC>q��Z�Ф�K�j�\�FOܱ}��X�}4Id�R��ٕx�@�{Fc��P�`��Wr&�u*̃�����&ܟ�1�I_�� ���Լ��J����*5p<��N�����}�$�h�v,\������mY@�{2��њ��縮ĄI7]��m���2grB�LՆ�̶��J�a�'�jscN�ܑ����w�3�Z�P��J��a[yi{���d15��|�4Z
�K�({q��8�^��v�ˏE�yE����@E��>��Q��9/����B9,�Z�� 1i�����=�>A��'�`:���Ʊ��µ��+�5*n���D�!w�� ��.H�B�L���6��.����@Nm�D���A�v.]&�����H����2�b��ϑ��3���)s˵��]=���fa����9�"��HL�G�g]���Ȑ�|�~(���K�x@/N�����_��-��cfzBx����8���@��nGE�!ܱ�4bg�ې��Sx�dn�1J��������|G �����;�N��&2^_Z���VtS�Xc���k2����VcH� �_����Xw�"�	�˚ɜUL�H�z4�LS1F��l�����gx8c�.�0�ʽ�����MV��ALS��q5(��iT�T�N��-�����-��k�U�_��{Y��ЯpG{?��iʀ��p�@�5�W���?����Y���}/2�aj#�r3ΩV��a��F����-�ݞ�bxt��*�� A<�q4S"�I�q-I驉��P�����9uoT�.]�a� ���%k����y����1r��k�
*���r�X��n������p���%Q�i6�`�n&�iBd���>2sJ�:�/��zɐŖ��۫�6}�0e�*��O��#��\��G����>%)E��+h���	i2�:��Ϩ�H�w6t��/^���_��0rO4j�m@�efw����c�|�M�e�k�Dq�WW�CR�\��K��4}�b]p~��0,�
]��֋�~��HC`�8x^�qG�~$uA�UQ��?��V���Qji�hoS��N�[��S�{��n�ە�_aݽ*� �^�/�x�4X A}�1�׻r�	��v~ϡ�:����1��d��`R�8�:(`��ऀx~Y��0ڲ�tBEϸG*�[������Q[zC��B7�w�5id�^���b�g9+A^�"�U��ȃ��$C�N�B�'��@�'tM_�%ǋT�m����ܨ(�z;
��%Y�,E��)\����x�Ž|�ۜuU'�C�;0�ɺ���Q��,��"g;��P���h����s���������ǵ'��
��iH3g8,6��j��Ņ��]�[����p ��#C;p��iU��ɛ�������Y���l�����i��!1��F:^ү .:7:�N���V���O�K@�6���|���������j4hJ�w���FCloȩ|�Cݿ�:�~��g�;�������B�t<��$��oEJ�斐��Z�[�����b�����+0�1�A�*�sWl�:��c4v�ۚ`ʺ�,iI��S����F�pt)A����jhP�4Q��WґE,c
P*]���>/��N��X�3��Y�ŀ��L�m�#�mO�d@BTd(�ߪ�C�T`N��5S�C<��I&b ��Yv���S�����}�y7�_Eؤ���E��Q��UJ���D�宇�OZ��ox��Bi�V���M�C\,P���y�JX,-�0��nR'�Su)��;'���#̀^L�
��/�^[���B�l��6������ J4�x_�z}w�UD�������l�[ڣ�E�I�4�Nq�M���;_���P���R��E)[��ND>BOJ_����c
x�4ؑ6�:<�a�ޖ�Sf�o��$d[�B���̾٦7��Jٷ;ˏ��P���gnI�.,���ķ�%.2�G ����ޔ Q���p�V@~�6�j{���E�6�f��� ���=7Xa��e��<�?���,���F�E�l��'��j�f�j��A����:�[��i$���I���J	
���;�z���A��z�3^��1�k[E��,��Zd��H,]"��	�8-a\li�XbB���P Lp|�����W�6�Oz��ҟ+��͚M�g�v}�ǝ���W$���G�|��ˊ�n���{dk:x\���Y�� ���n#4�&����϶�Q&g>,�0��V�gzsD�J�����؀np^�C
v��6^<I�y��Oy7sZ�[t�ܸK�N�gxB��Z�>CЩO��	�W����8I�*'������h����8��/W�|W�K�*�l2ϣzĘR���	9H�}�H�WC�:�����v�[���E�M��4�8���0�Pݾ���i^�tZ>Lէ������n�yR�( ����8������cw�{0��Y���nc@�UKI�#�7�N�.�f���ө�\��֠8���o�|�Ŧ��v���Ʈ��j�:�W������s��(q����:Z��:��B~F,S��'U<�����R�k����n�ζ���M���x`J*C�<{�uL�O�G�)�E=t���~o��9�Yi���z�>������C]����/��.Cl ��A)�
���RU���pN
���:����+:�n�k�cg�AZ�<�oHrQ	��(�؞-�տ}s���$�L�N`k���nM�[�z��'��S��n��;�~��c�o�&�&�3���`տ��5���b8�rb�3���]C�Վei�Q�Qwj-c����������g�T�,p{+���-��2hzو�7Ey�6����GuMw��� �y3YS����oU�/;\['�����������d��|�I��V�iLH�*�k��Փł��e+�u��*j�0�ߒ9��[�ℑ�T�����(#��9���:������O͝��T"���;(
f�0���O��8����Ю��~� ��o�I�m�å>k���w�}K���M]��`��&�����s��+�sB����\���|wV���[ѽlgH�&����m6 ���Z�⥋9Cu��
W�PWh��hqS����~+p�
��t��X������<�i�:$�1�j��k������0�'� �g\qb�G���Ty�����)<���ko�d��v/�A�0�B�ڕV!�G�I����4���$�J�Y"�
ݞ5����G .n�@
���hL*���ՈL`��z��A���{���"#u�A���2�,v�,�3D,PtQ:.�e�p�;}��ݍgQM*��K�3f6���� �� T�A)Hs�h�`XSi��OS�0�,�*>+����o�5��<�E�~O<��_4DЩdI/V��!#2|���K�B9!'B<'�x��:.��[{�3�;v͎���9or���ͺ�S4L���B3��2.�q$+�B?He\�����&�5kǞ�[G��+��.�T�<���Y��"� �#��B��y��G�`�V��j��f�3q(~}1	g�6�u�i/�'�ǅp�UT��Xs��Q��ت�
-L�6���s��Z�v��` ����w��� L�Sq�x/ko��=j}�:_��M���j\�9n����ˬp�.�iėw�{������䉣�`ȃ�
[��=�矍z<�ʟ��ˤ��@�fjO̷(��u�~��5�%�B�:�	�s�~L8O4�a^�]�o�ْ�����5��=f�j�<.�0����t���*�1����g�F��.F�$n2O-m_�i�Њ�\51�D$|���.R�R���4Y\�P�:�
'���"�]�dOV)��^�p e�iz�%g�?�
��Q1b=�Vt��?���|Q�EVvU;�~k�f�qf���8.c�¹ ���f��\a�d��2[S������e躉���X&J�h8岉THxb�Q��./&��hCs1�U,F}ͤ�$�c�/�%���bZމt��B��-U���2��֑Κ��e�����/�@�@�g�azC\��c�!����?��P��_e���.jf�a9��m)�j���y�Z~L���5�hv�.Tz$�&Zd�'@���Pm��H����%�|�j�d��y�z=n�
�@��X��2���Jh ���ɡ��I��j-����dcc㩎 �aB��c6O�"z��^K1ߤ��T�u�鑈L�T¯�phCB�[?�	V:U�R݉}V�����-�)��Xd�y2T��1l��YϾZ���J�3`��5p	_�FΜ��7����k�+eѥ�+ WD��(?�m��\jq����?�a�.��4�ū�a��������П(��c�w��/��RTѾ�m�H�<�"=�7�0�mne̠^ ��rn΀!�a#6�}M�$K��㒽N�C�)�O��Xz���Y[��j��\����iҔ�y	4EV��t� V�J�3>�����7���k[7cx:�l�#���?��/J��Q�ZH=�L���kk�Ѷ?��e����q�춅p�\�l*�d�����1(4[l��1��q[ui^���W��?����@-�c���˔�"k��-yo,���-zU���`V%g���Vn�;�KC� X�+�:�8	\St�ӶL�XEC�a)c
�����`�ʊ=��_���� ����vB�t��>p�b���G�gr�ہa�͝�������퓱�|F��s볟�>@��xW�:��)�����	f��Z���_��'&�"�4��
�m��!�v�&�e��:}�g�H��Bd���0T�[�>�@�O�nXv�4���	�ĝF��?܏A��	��0����QB��R/2��2��Mfȟʼ$��:-/��S㜣����o���{�3��c0�X��b��]�K�[ok
k��9zH~�n���an���	#�^ﭸ.�$�5K���F�����n;F��s�P���Ӓ�[k��}�����+�~T7��%7�UI�쑅$|qA�:>Wj��#zV夌=Xh�V��dnr7PFx~{���4�n��hi S�����R@u��}w�_3�S�ɿ�08���r�u6g��V"�άex�Y�لs�.�<3�"Ѓ�5����/��IKT9�T5ζU�)U�D-�H@�f�Qݸ�Qa�3!� D02�4K��]��h��J-��oup��"	�z�2�cD��g����@I���bw�y��.�[��z]yU0���_2���B������^�]S�ٯ���B�B�;iW�j���N�1��Y�^��T�[~F"Jvq@�ى;M��`�����n�0�Rϐ�'�IJ�
�����O�����خ�Z���~ڑ޿U�N����U,�N�r����ڷ���I�e�S|P&������B�������.E�Ot��}�wR�z��b�M�i��h���)"�fD-?"�N�n�o|� �5eP�!��im#w'ڛ�~�ֶ���)l4�	�����]F�_U��|��e�=}e��^%б}+�yñ����B6�n&�砲��<5��#�].Eo�t���7������:�:�c֦��e�j��I��x,�����Cb��¯p v�t@��,g���
���B��&*�%�ﮃ;�11��I��'w�~M�)��$SV>4ӽ�z��*�L	Q~�*%�0X�Sz}�X�����PEbŉtG=�0e�Pj4�5��J�,+<c��7�����z�8�V<�u�1{_3%�-�������ho�8@��bev	0�Y�L;� G�����8`M!�����a׮����a\�[���}�t��ߔp�B^��|���z!y<Z�}i7�| L�:b��L'�}�')ī�:g�,h8���{Â�if��JnWYE�/W\�_�Q�7~�`g�U}�ki�p�*�ޏ,�q���{	}��z��0
`�\���^G�@�@�_���̣A����ǽΜ�e��>Cvg�D���Q+�#R�8P�,{]Ѝ��⇠ ���h�[�E���n�*�yZ@�	��EL}�����R�����뙀�8���A`���o\o1�թ7��~<7����X�M6G
'����>[�����ܽ�'�����c-�����'Δv��QA9��Hz�g=�T��0��? ��&:(w˺�ӑ����3�]j�?*�ηk4�c�q�K�[Q��'�Yo5^z^Xܾ��!����+&��_�z��	��6
�E�~����?G~+���±+4|;��Fd+�8�x�����	���������,�!��<|�[7���KF���h��M/�Z.t��#��얽�a`
V�"��� ELzWN'�b!��3�ɴ>��SF����]v�L������w��t|�$߆��Ɏ'�e&��pd�Bp�`e!���B��z9;���z|��i�8�zx���g�w�	�!�����	/�M�^��Xs���Ƌ��W��rȖaC`)^WE��v�%?f��Wx�~������EXk$L�Q8�#l� `����ܗԡ'���_^I�@0��ތ��(?�hn�LXiw����R>� b�����2�h?ޏw�o�Е�pE!�se�	����ٱA�#��a "[��vvm��䜉�PbQ��).�&Cm)��%t�Q��� 	c.R����S-�v�^���y�)�g��RV�9�W�f"�����)O� �W��|��t��*��2��+����Q�	)�9�`��N�TOܟK��m��Z��E��'P��$NP�ɂ�XOn2�^��悆�<�-�.�6<f�̗W�z/^n�yO5k�K�=�˱n��DW�� ��1�J�UV�S�0Nt��Aʷp.V�5b�J�{yj�K֖>�ٓ>��Чf��Lb�Ha�k&����x��%�w��So`��<�����R��s�a�䗵�F�[��9[s�v?�!ʛ�@7�O�����_XDJ�o��u�):Ǣ�:=�<XH����g��X��D�ߠ�7���W>#5*��G���Rx��$��p$uh�	7�)��y1��ߑ�i��}��l�h�A$d�1�,�����RGп2>�1��c���%X��(�P�!%&�N�Z>d=}�/	je��+��K�/S��sܾ�@,Q	9y6;B"w���E���o�:����d{4��	�>���/CGd7�4������d�S�#܌��F�(SڅK����%��Ԣ $�hrV�p�X����]���J*E<�I��e�����;W�!1���k�)����a�9��R��'i�|;*!y��R�1��s\pg��B�X?Q��^䭥n	�����eq���UOC�����q��4a	�o���,�Q8��B�Fɽ:_�[x*��d���[�cʏ>�����1^~i� �Y}�G� ����c�/
����P/1�Q)i���Y�@�b�pA�0��y�m��Yud�l� �#E�J�CR�M�#(� )r�iL ~������%aa���7�ńFጃ����M������o��
��W_�� 7-�ț*:�M���V��F��@���W��?�U�Iyš�Z:]՗���8�Dh���R�v�����H)=N��
��O~,�PJNzJ�d��6��M�:�n�BQ�T��x@tZhg�jR�j�B)8�!�M�KR����3
o����1��tfY�5E~�˴��p<	�]�E/�a-xy>P�'{{ �<
L	�#t=�Q�����?էbJɘ̝v�ZS��1e�9��Za�g��K�BR7|̽Y�S�ꤥfǨ�w�C��J!Da���@�1R�gpby��dR���9e��§�̮U�D��q��e�|�f�K4	�QӘqa�.��`�"�'k��w�j>"; �4�F��Pp0�D��rR�-V�ME: H��ӌ���R����|�y4����'��8��!��[!���=��A%\��@�.�6�[�Y,��8p�u���K`7�_�B`�7��;.�Z�'+{��������nu�h1�x�VK�*�յ����1zN<s%�d�<�w ���a<`r� �|8@���BW�g�ҭ�m9��h���l1I>��:+��H<��G����[�4�$���S�ī<�I��6s@x�&B�fu�`�w7�Y�J�1g��<���d�X����4������wɦ:���b}`c�.���2^&�e��?R�'օA����7�I_ ��5۟���0�^���`7Ԏ.���-�1�r�%�5���2�������+o�
C�`D�r�	5�x��&��Tm���ܟi�Nx<	S������%�^�N�:�|�7��3���^�r���V
��!�Xn�;+cU8Z�)���D*aa����"]���?:��|��܅��e��^�k:CLR7j�1�y���#",��=�>��& ���`��=8��8��	&��h��gտ��Zлϲ�Y���X�M��Z�֑�m�[m�>d�<>U���&��_"�!`��݃Â(�}������B��A�,"�x����-�\���O�cv+ɦ�Q����
 ^˸B&g�ߤ-|/K�re��+TP[����LI"J�oQ�6llL+�FeA��`�9r�>��ۭƥ�{FtC^�f��XF�B7/�qت;�z�l\��/�����(_����p�J����BA������yI�O���`&��#v[7N�.���uVEH�>oj4(:��W�"����d��h�[޽�>��4g��3�=/���RM�L�^qk�@�n�2��=�:O��^�y�>V����D�>~�I���1Gd]�&�rdhF،0��Ka�����/H�Q�_7�O� ꘚ��U1���.����p��߄�����"-u�oGZ�P~�TC�K��x��M�qU��9�7�\�vm=ǅg�b]ѭv�e���9���%��<e�3��Մs�@���D���� U���G&ܷ�m���50^�{��2�ә	3Q���|��E2�U�w���.��rB����Mux�J�E��x(�F���d=5�p��8�����RCY��2w�|�؀������>v|2A��Im�uuM�L�������[�>5^D��hR=6�9�m���U��]�`�@ '���ɿ�#�k 4������0��Z�:��3�^�6�>��qoZ���j�������h_��������������c|�G���e�N�.��,�ڇ��=v:�ʃ��n�[����nڕ�MY_��\rj�x���o�A����wg�F"�Z������jZ�����ޟ������i^��&�G�Ѧ���j�:��6m�h0���{S�@3{�r]f~$�<]p�Ơ�����E�{�8c�_�U�I2�+t�#�'ˏ���2��`��ǌ\�ۥi}�Xg��qR�����R��I���
��l-�M�Kk� M^��\�_8����ɢ�>���DMH�E��z�F��1�r� C���M��٭#���YJ�Rm�a��0�z/������}�@�a�� P�B���}T-�]=3I.��������U��(��/z��G������w��5�KHx�C0�����;/��X}�-gc�6i�8x��[?\������!f����fB�i�^xėm�~o[�Љ�	<6������y����o4&�Ҝ��:m�R���DS���х�ӥ(������������
���:h����yz��P���1	�r�b��a�QklD��ƗX��Q�I][n���C|
���6-���j,�B��_�N���<K�i.*����I���1C��2��m�YA���+��2Y�z%<�Br���Uͱ�}	_�	T�Qz	���}�@Z��"k�tH�2Q�3L��(��m��É�ȁJ���S�e����ogwۃ�\����5U�!v���^UG����`�8#�<#�*Q݃j�&Y+J��ՊbZ3����<��_�WȈ�F(���[���)c!��+�%_V.=m9���	��v�z#��4�J���gU��d��gШ�&Gzh�aiҌ��$/F���Zl����i�H���TZ���B��twjKRu�D��	��E|�פa4]Ҧ�z�������@jy�����)�j���G���Ɛ�X|�M�V���mq�
�3�����a�����4�$��(u�g�A�b>��x\�ê���!|W�+2��Q��-{s��Q;$H�`�Ǜ��	��%�Â8cH�6�~���b���q���i��Z�g(8����y��Mo۔�C���NR��D!����F!S��9���p�)6ܟ\b]��}�-K$���<ֽ�4f��^��ߕ-���=�΂�]\;�]�U�Q��YI��޶��-q�0$l
�Z�)*�� �%[��C����S �T�ae�J��9g�����f_^yvT%���E��*_���߻*Q���{���)�D�${N"0|3&G�!�f6k�W�����;��Z����7��[I��'�ƽD�}Y��U�a9�#t_����,Io	�FĿ���ĵG'������k��B�����~h���
	�>fY�Hs�q@G��x�ـ�=�[�;h�X���1��� ��w�L�&��0/-�xxg��Yؗ�cd�4OA�G��Yq��8��&��%-��T�ҫcX�g�]8i�H��J)�no3W���'��܇`/=�˞�@��j&%�:ʈ��Y�vN+y�{v�>�>J6dE�>5�I9<]Ԧ[N�=�L��36q���z�+}�j��aM��+��i���{D �����qn��еl�~0Ҿ>׵�y�hB�y��ix��:Xg�\���R�_!��pS��k ��n�T]�H�	�%���ˑ3ì��T61��U���Q$�R�*��S.SG�g8|�3ʍ޾I�a��$e��P='p��!�-�Ο�P�}��Z����:�S
W��8֍�8��QvƦ;�Yi�h�]�@>�+��)�.P�]W'X���eF� C���<C�03�����$��j��.��lq	<xb0��Ԣꨙ\%�ϰ�^'*���;����(�_"ԼCbӅ��O���|q|8u�Uk@��i=e���J�>��7?������v�٘RP��Y�yV��)�]�T�َ�rو�֫�k�a����5�V|��FZFu����o{�0��(�PZP�lS(���o�O9О�n2�H�<�W��2�r��2����2��C���r��oF�F���1?O�e���\^���̅�5��F�~Ik�o,,�ʈaVF){
S�a�F!����f}p�s���@&��9\C�����n��եm�D�EȧC�Q�'0�sH�n{�l�S�ք�����zظ�#o���+�%`�ģ,T�]:�Y]\l�V��
���s���m�ao��M����S��⍓� <ؖ�;��-�]����B^W W;�*|�:��#	�9��s��/%q=�cÈG�)Hsp�����Qq����
���
bk�X�:�yW�����u��*�zKA�Іǁʥ���M���g�2%j-X��%d�4�Z�,mDo)���v�s⳪u�"N��I!�n�<��K�39j,��1S���}�(�'�f�j�@�	�:Ԃ����Jy��<�܆�Byt+�`�����
F �4o�c��.68	�kk�g4|����ٴ<��g�d�B�l�v��'b��v���4^�I�"x�\|��5v�=`Bڟ;��7��¼�]_����SR��$�`1Jn��e�²�/�9m���t��"�����a7$�Qf�>��$+�W�#�?ݬe9rJ�/�M�h����$��z����L!>n���є�����M��@�k���g�ݧ6�2����$E���o���MG��;TL�����x�FN1�/��}w��J�,s��=�R0U���߼J��kmu�т ��ճw�� �N�`϶.�8�d�R�><�im��઒O{N���g�z`�(�B�,�u��Y��J�w�R�Q!�Z�J-a��4X�5����D;� �7����e�1����Ǣƌ�^<~#_����R���P{J����`�Z�Yx�䝨h���W����!����I�QY�˸���j	��(+������=��pz!�Uy���^Yv�gC���X���ɨ�x��+z�0TZur���t��!X�wҒ�3���܆?��ӕ[Q�9�-���I����V!�#;AV�۠�� ���[ّ��N����"L��^���ΞP�
L��1�� ����&��XH{{Mis���F�u����SR/�H5*��G!ݴ�j�����9Ƣ��61��~7Gަ�fOXNbnV��?�1T��:>X���	��)�nIS�,�����#s��\>5HVrL6Q��a�@y3no��4Lj�w��c�|Z�
B���&����d�&�)�f�_�'h����M]�-��CC�8UO���Ty�i���[��a���������!ĳ��Ϥ�Uٞ���d�u���|݀�� ����.���mM�*�2'.'���J?6�tp�}���1�\t�	knO����0p �|v��o��!�!�^V�t/��I�|��M��P�u:Uў`���dv�tx�?+����<��=Sc=�3�Q ��wh�ѣN�a�v4C���*�+>B&|�����D�1bg��;�'�~1cQ�B�{m	�4(���ڏ}��a�����ø��X2gc���`�l8 ���9d<O��$dx�NEG��'���n1�"뢀�.���DU�K�KJ �����B�8_��$B�`�M�
�������F�fë1�|$ؘ�KJ���@����{�I񺹬,m?bC���9�C7�؍h�)��� 6��}���'�cf?�\�2�/�x.%r��/*kZ�=S5�����Vq�Q�s����MҼgQޥ�N�vslt�\+��(�,�w8�a��,ɬ!t�6�
v�����*H�G���t��>�P��7=N8��M�̘h�^�r՘Li<�W��̡�68�%�����O�k����/Ľ��u�+�cJd�+�<�[Hn���R����ʟ��fkli����q���m
!
~�M)Tj��`�k�#5c��+�z#r%�m��p��|�\�a�&��#�H�ّbD���*��7���2"�������·��w3a�4E����w�DE:���0Zi�9�й��d���Xk )b�8i��!��]��޴j��`��$�nD�����
AB8��A�CLj����ѐ����� �`��	����̛��`A �K�r�.��v�����!#�pu��t���u���d�H���Y��=�.�B��XJ��D́Y=_�5Rn����*_���������[�	Z� �K>B���y��m9�Y�e��2�1���l�D������?��]V��S "S��Z��6cv/V#S|[�ߴD�����w��9=&r+ţIR�	6ȶ[�o�Ϗ�p�D���N�Wďޕ�%�uH�P}��� ���z6\�0&�2��j�Vr$����������3J�/�	�NKG�<^I�\�Ã�"\É�
;XJ,Y���Dw94��Vo�v��-z��<��ԕ����}Tv����.S���M�27|���9�]��������L
���IČ[����?�q/�G���D*_ꑯ�L4O�F���[b���qx˜���lo�ͤI���ѥt(���ݣ�y��͂�u�7$fw�v��Q�O�7D/�c�f�H�L����������Ʊo���2[�+?����j�l��!�yY
~��=����M��N��b�_��3a2�o�-�`9�W��E�)�9��_����c�W�ll<�Kni����O���
y2X��,�R��	{ܳ��M5�Ì5��ɼ������T`������Q?2�J<�&�ƹ Tȑ�����?�V@��XAlX{��ڔ%R�n�;�k�Oϣ�Z�THX�*k��M�UY�X�?Up��Q�e��u%��?�Z���K���'xr���^�Y��Zjz�-J�Ь~����k��Js��
�,{Hzr!�5_;y�ǚ*}���c���R,Tx�s=��`�������)��DM7=�-P��>�!��D���<W���ɇƖ�Mv�d'�:���^�;"eE@��BbA'#k��t��N��+��vO;�S4�>3��_0�����O��YQîv@�nm[�Io� �Ƣ��
���iwn�Y�	��Wc�|�B�6�D.���y^�(�`"�V�Ӧ*4���	ř�5݋H#j����Ɲ������:P�?�\��iH�<�pϿ�h6-
�N��/9TST��rmO�	ɍ�Z��2_��%{Z�ߨ,���a��fl��$}%�f6ȯ$�T��dzd�n����V��I�kBG��c��V�a;"z���~�ب�k�d�� OO:���M���ͲUl�J�b轖WkE���aH��ͥ4��̆�KK�GQY�:A��	����&��;��F������	~NR�n��Q�y��t*�}"��2_��{=��K��8|���
mj�W��m�����B�u~q�1�h�a�9����3~(M[4?��(��@Z3���ެ}-5��Hɉ������"�UW�n������)O�����{���%�AhG��?n8���""�Gm ҂�Ԗ}�Ǣ@��s6�i�ݠ��q�؏�L�]S�E�mӹ�Y�Ϋ��&:r1��A�Ƽ/��,+c=��Y�Y�|������G_�8_��@�Di��_T^��N���{���E�0�C�刪uy�)}�ȳ�%'��bOC��xk�9�Z�k�+c�|s6��ų�����<�]�!7�3
�߳��m�nyy�F���[ݖ)���xp!U�)-q#�eޜ�A�>��K�w�V���p�Kk������<�7�+Z��IV`L<��� '�1X2�n���Pu�3���<�D�al�|
oa��_��]��dK�h� O����Z��ρS��Q���UŌ�����=�Jc[?��x�����LXߒ~z8��#� ��?Z:�ì� �צ���ǃZ�O~�7<s^���-2����v
玥GɃ������4���/B�5����#na��
�u�S�U��i?�|����[ԋ¬{/~��s:d~:Y;Â��6�L��%Rψ��B�A�F	��6�' ����H���s������e���~�f)�a��E��C�Il��X~�ӵ�^<cnר���fl����6�L*M$�7�Of�����|�8�e�ߊ��}'<��{
�2}m#�����0�G�;���mV}���z�s����t�e������wb��K�Z=y��;�2�oZ^"�(�YԗܧAɆ�b�o�#�v�x�bH0NA���Mӛ��?'Y'�e*���7��u�؃4����3���#���6��oB�́��Qރm���pS������1m�|���S]�l�U��.���Ι�; ���g�D��X,�蟫"B�|��n&�'W�j@��Q��}�;����յ���`��Q	d'����<�h�շq�����L��y�=p�>�H
h�ߌ4y�9�"��j3J�/`�v�ft:{����Tg'#׋'�V��a�FS��u�|lT�깼1��?ǭ���V�ԅ�{d��S�,��� 	n�p?O��x:���������z������&.��KA��M�u5�		7��s�^�d?�/b�QPh��e�|�Rx��8��G-T����]_��og�������E4�	$xp�#K�戉�����ς��@�l��V��y]r(�/BY�8cY�V�R;5�P�@4���ћ��ԯ��z�z�K Cmy�'n���E'��Y�_��ؙ��S�j�\�4���(]�� ��p�G��H�G&�Y9�c��R�Cl}�%L^��2s��6�0���VwC>)m��/���35Aw[�u�P�7v�R��UW쒷��t�|��
yB��B�UK�zFZLv�ܝ{�
;�!�����K��A����䍑�R�b�!���ȩ9�[h �;F��P1����UK=�@J���-~�t��W`
~Ŝ�[�(�b��Wc|�"��O0x��h���Hu(��,H�	ޗxSv/%9�ǲ����k���K�2�����#�E�{�P���7�pHlշʸѬ�ޫ�@R���%#��t�ތ�CGa׾�T����b����ET��W/�	s�WE6C�F洇�g�n���l��"�HD~�Q��0��\�P�H�/�B���E��������jI�?��3�hef9�������Ҁ'������u-i]Z������8xڪ/Օ�2����wb���#k΁44��N�I��fA�f�����>/�)ڥv�B��������}�U����n�YE^����w��CӖtx����8�u�� �o�2���`|9������*�o�6|�M��4TJ >��-�^ױ�b:@���J����_��q�$�5Z�E�b�/��|�0���;Ph��
���R��1���GU+��)�e��8�l�`ϑZQw_��i?m���3�5ո^A �~�fÞ�����*z�>7ޟ@@�d�I���f�_g!�?��,��m�̵���C��7yJ��'��������X)^z����rD.��n� �ʙ�v�XSG�\j'�'0)�.��Ϗ�O�dq�����2��	�w���СUK�!:����Ų�Z�P�!3[���@�=��.̅������pq[9MJvUi	�	��bYi=��W�\_�2k� �ߘ���{�Ւ�ln{ތo��6-�֝�H��;�]3؎6=yg��I~FAdVU���k/�n;�>�i#�YP7��0�Y����!	���W�
���T;P������]UV�y���뇖�28�9<�WZ%l�%��d�a���$�rHL�'Yb_�;���`�������Yӭɽu�Hv&^��l�<�C�-<��SFz]<ϊ��q�ྐ;c(�\�>��֦�#9�T�˰ɰ������Y+V�y��a�$��>W��WP��e$2؟�����t���/�&���(Q�S��$�-i_��"�-k�(v���k�?���
�UY���,�`V#���1���x�2㱯=�S�)�O�1@s�d{2>�%S���#�.�?0<��#�ǭ�����z��'; y�zj�Ȃ�w��o�apW�ݑ���5�n>�{
vx��/9�W�\��_L�3�M�-#1�P��H.���W��i.�kΕ3�!	
Cl�y��`!6�-���O�N��7��1�R��3���#XMDT�(�y�[0���50-���y�z�ӫ{�U(�F1t��iePm[���*��>���]�B�L4ē  F���[�p�a M.+r�HvEV�_�PTk� �B�G'06�������W6X�54@����A�]�bO�T<��Ud-w�ZX�A�K��	�� "��b���X�����T�v{+�u�.����:�A<m[U����0�����i��zF���w��8&��)��O�'Su��̾(�����A��b0�[Ś��\�m�_T�o�Mk��aV�M?�.��R	!7i�P���
Kc��	|o#6��)���� 8o\N���N��<|��|�hƋ뾋8w�ۃ�7��b�7�_O�ӓ\�����~M�ZlC��b+a��e���/��<��|e�4W~����6d�Y{⒓�~�B�
�n����m�c��Y�V"^v]�����l�y��z��&�嬠��8�Q��J��M�G����������>Y�R4��[�T�kmxGf٘�	)�ɜ�9 ���
���Ӫ�}��D[���4YiJSb,ND��5Pzo��Z�~��)��ɯ���t�D�����y�r�qۚ-���N��ȕV��FUq?�|�b��N�:��H�T� ��2��Tn*��P�����o0IȪ<-��$_J|M/�MrRr�j�բ��2e܍�y����
I �.��!������w� D���0�/h���tr�[x,t�}���<H��,]E�m�4>��Kb>�<�_ ;Ԡ�.�-��_�˖�G/p���ȼ���EE�a�W��ih5m(�X��<�p��=�"k�c��X�IP��0|4A>�9���Q��J�&֬�t�	�fԨ��f<��yz93b��*s��2!�'B�ZR�[�����	�t��T�P]: *��rx�l�<�s��M�鬄9��4�nX���W��R7��l�o�����xǻLA��JA�����Q�1m�R�	�8�TށZ�Ru�ν�1�34bb��+;9�nfh:^��i32$ܒ��������AZV�:(Q����i��׏��W��i�����;GG��&���U��>����r�K��>���٦kQ�3ܼ�����w��G��+�/�����e�����
X�}� :��[��������6��Ԗ�$�uI������ӽ��hр�ם�DC��:gH��OT���?��.0;�@(��7����B	m�P���� S�Gm��H���	���n'1&s6��������_(c7Ž%�g�Qx��^P(�G���5��Hsx8�����R;9<ʐ��5���n�����N�,�ޛ�'�f :�,��X�!�K&�M�$ ����?�`2��L`��4���N0�x�0���DfX]�v(�H	��w��&�p�!�f8��&�, ,Kmشi8����ҧ�]�L��=
�_���Qn�~��w�����ft�R.r_vj1|w���@
|��혊��u����N(�JzĐ�a��ʤB��L"�ץ���<�J)q�e��f���0r��7%�@R7�R�"yUyK%Z���\� 6{�gE�o���%`m��zODg�Co�`5�5/ǅ���+���+P����L"�%�G}N�!$��Uwz�����_�&?B���w�a��u����1�!��fwO��{�u�W?��y�m�u�{� �b���8Đ::�~�q�*�lp��&��,W3+��&���{�ɶF?�>3�֌>�t(R��ޝ�>4�!7���mA4d`�\Opp
 ##�_������rom.ܑ��lT��}j������U����*5�?f�ʸ<��Y�AT����}�#1�ɊK[kB:p�U9�[��q�dMEFhL����=��Fͪ})���Y�L�&�h&0�w��A����$�z�ɐ�d�S���xC�������z��4	�D�ŕ3�]�N�'Ǉ�&��<�u��4�[7(�[�P�5���>q��]��R[����	u�����?$Ʒ �Ǩ�1��y~�S���y�*RD�&��X�~��'���N%��yVݞh?,���*�5�y�АR�Tӝ	]�GF�|���ב�Y��e���ŭ��b�S�}�n����6(���,f�pb�O'x;���ð�8���B��m�쒋��d�[E�2'9�k�^�����5�T���M̥nIѪ;���I�5�#�9ba�{�b��b�����6�ރK	�K���!+)@Nd�"Y�[���.D���{̉��ˤ+���#U�{�eW��G�kk�x�r��m[4۴(� �'��`�5��+2���l����[��u�m1[��I�ye�6N��73�b�7��W���s�� ���DB\�ј+─���⎗ѷ�lQhx�CFn�t�c�bW��e#a,.�$��YWZb���N9����J�/p#^�M!�b
��Z��.4��ga�i����ܝ��@�O$kC�J�(��|�p6w�b�V�e*���d��U�E�&A�NMka��W
�$��;�h�?�~x��掿���ݩ�l^��j� F\.���t���Z��W>LΜIPxb�<��L[P<����Z�vWY��YW e.$S���v�����RAW�+t-3�ײ�ARѰ{؂�9Ϯ�����e7����
U�<T0|v��'
\S˛��v���"x�I�Եi����ʙL[�Y˗��j�2ge�qL} �1�f�&L�L�.�*���;ԎĨ���N�dy����.Y�/��c􌟥�Ś���jiT��ax�+�e��@Q����~�nF#W�4�s�?	0c��t���-I��Q�]�]�
͙ ���&$�;��w�|dQ�66=��zzm?L������831������skh=`�終g��)���t�o�a��_i�õu:�k��LE̋Yr�+z@�6��|��:��D#�)F�|�N���Q�b��b|Dոa�r �G�oԖ퐳_�)�LEJ�{���ט�4{�y.����t�ƪu�����9c��o���B�x�m�MkomX+B��G�	�m���͎T@���p��2A�/�D�ͬ�Y�\�=zl��(Ŕo1�(��щ�O�g2����ϓ)csM�<�GV�\|3|�z�{6c�;�Wmϼ�(x��w�2[�,ASn����� <ɤ>�{��t���jCK��Z�3�_f?~:�@��|������D`�5a�_|MEA?2�M�?d2̨��I�c��b}Ǭ�OǉQ��>,��6�;�K�H�h�G	�U��� 1�z�b43��Z�s�i:׫�B�8}�����׳u��R�1J
R�V��z��󢏓pcH�$�O�o1��rD��$Yd��l��g�^�,$A�G���(�F a��������}�;��R��h�:7�6Bwe	��?�<nvܖ��(0�v~��6G�<�������]^�mւw��ވ�o�p��'נWx�}%��AJ%w-�+��b�QR�nN��pE^��93e����C�"��o��K@?H^p^w}��f��V�Ro0�:�w�Jt1¨��n�@6�a��:�}q�MHp1��N�︴U�zXN�v��q����]�&�r���%��g�a|3�����L����-6f�A�m���<A��ޅ�#Ζ-O�_�b�9w���o��'o�C��㡈 �BJ�ލ"��Vp��|����U+k�[̽�N)��k�t�_��s�sb���T���������� J���KB�ؓ�+0�^Ӥ�?3����٥)�7��e�m;cj�A�1�@�#�ͅ�mg���8'��p1�-���z턂�}���!����h��
�=a���7�1 ���I��u���2������������|�V�IA��[(��<�����A���h��;m��'G�V_�wd�~�D�4t�%���z��ɮo������6�����~z��;�����Iݜ�:,f$�x�<�a�qU��#t�����H������ȉ��}�v|\�-bI�3��'��f|S�	��S4ط��9���o�uE���	�Й"C�H
�g̕U>6�L�a�1D��Ε�-�5F�솲5﷣�BGhP��;�B�?}�z3 i�C�az�
��K$�P�R��8��"��r�-a>�͝��>�sf�~�Q$'	0<���'Q�0UV*�U� �q���ɽ'��+W�w�8���ώd\7��]T�z�l������T�|IC-Y��G�ܘ ��u���S��Ѳ݂��x�����M����ݨ���q�m�U�="~%g��Gt�N�ٌ	y�~�t'���$���"ɒ^]�����FX�f����НL-��|"�@�!`Ř��A�n	�_*��"�{�?�2j�hj��mh#d�`�����$!J5��>jb�]�'l�*��x���+I�'�]T��d�.��&f)V�co��{�O6:�=8�O��Rϊϋ����\h3I;��x���뚕�E���xݹ�+�7^2��	��^U���D�4����t)n�UI��U���w_��\uuֵ���'�C��D,�,71+�Һ�r���O��u<�`h�\�R!�rh"��2��­�F���xb�,�?K��4N�"S�k�-�,r+�`=��!c�(��k�jÉu�<�X9ZI�0�BX��0mo|���h���M~��Qw�6�Un��z��HN�BA�g����M���wPs�����	~��T��W�]a��c��5��P��	
�Z��l�JD�P�cէ$����)ˮ��.2jv/�v�T0A��DG�~m�K�c���j�s���.�����R�ZE>��l`��ě`w� }o����4���	Jx	?�Lx��C�]v���'j�ع�L�����cҳ��	+|�#���Y+����� I�j��V���)��������C��+�?����!�����I�e�[��'�]"h�(�`n��G��&NԌ���SzLm�������+v��Cv�J>Ⴚ���<�ia�A��x��$FvdrO����2IvQ�����[�8%� ��T9���^�YR١�s������n8m�j3)-Y5�3O��8w$�J��Sr�Z[ǔ��Q��B��K�.�kB��/��&�#�������L��fz�-*�Y!��?Rn	�S�rX�3;� ^l�*�6��ZA�pQIdɷF�n�|?\���1~NǶF3r����h9g�f~�$��ê�q����lYG��E@�j!�| �}�p�D�,�F���y���u���Q
���  ���o�ϒ��sS�YPUY]��B��0V���nN���;�D�8y��c*@IR#u���XYFv�<�#�T1��|�� �b���)�$�_��e�<v�.s|�t�*��3g��η�DW���1>f��>�=�=TJ��f��zz_k����{�V�Ktz�-A�)�0�H�`7n�T^`��+틨���余�F&afZK{`R����ڱ�}o"�y�)��p�gg���_W}[����.�Dp�D��6���j���D%�I+�8}\�%ԬF�*�ur6,N%��R�F5lt����l% �e�����)C��xv@e�"I���_�d8�N�(k����T5P!�ؕ��B�%����@m��c {���6|WEG ���Ei�^J&Q�>��4r�h����eQi4��)V��U���h�i�Fv�V�p����L������k{ >�B��?A�y`�����B)P��傄-y�:O�������K���b����@�ٻ1�b�Yھ��<V�r��}��C.��P�^�H���[[�\J2�Coi��AS�L�$�c�O�N�����Ï�{�Ff}���O0�t�48ټT�^V.nOϳ3Y(���&{a�����c��P�l�(��|�ܽk�$�¥�X{�s�tG%����T1����P�3��PՑ��LIf	�rDs���|�pZ�W�P�)Ta7f�^zP�����!���Zm����E������mS�^��yed����C5	��ox [x�W�:���#��
�,���'�5=�f1Q3!+G�p��V����kv��c:aP�����K��D��:t߶������/K1W��Yz ���sf!3�ʰ�1�u0?,b����������{�uo0�¸��_�qP��j��,f;��_HI-4j4�2N�ޛ��Aw���Y_
��Ul9�U�ɵ�܁.(�|v9�BъlM�ǹa,$������"�=�"f�b�I&K^���:���2���3Ү��K�FM{�o��/rd��V��*젿%��H�H�+Zo�¼y1f�ʧ�����&��@�#����iп����ji|�2�X��|ed�'�P3��Y�����:�շ�V��wLӽ�������o(�,��UX���X�tc�T��J&)�^��ю�KufV)�n�#�Bq����eݘ�ტI]������}�������^����|G"���t*���M(�gN<���=�
�;���ǎ��E�NN�
!��$��t0�h��U��2�Ƈ~�qv[�~�c��zV�gJ�d=#�{aź���X�i��j������"��4>i�*~�{���~�^���{_s� XoY�@Xwa�/@h�$�"PyZ:�4�nuFi��/5N����S�߻��/CY�V�����㠙�ǀĐQm�L�mx��`Ѭ�C����ȿbA�Gr�.+x������tS��|m���0�ܟ�x�2lL�Dԫ�B��24����x�Ξ����B$D�O�8������(T=�[
�g8���F�n�X3���6�[��?���Ҙ�2��	"���.@�%��a�-�� t�Zh�!Ƈ3��K ?+�;�4\��X j��_M4���T��-.'o������\�ٛ����x����Ӑ���O0~4�*����4l��G\~ �9A�h༂X��KIo���u߾���-���M�Jo���fI1��,d��z�j��%���4�ܖ���ơDSg|�5aGd]�}��S��>N@_ޮs�e��[���}��\���	X�ad�y�����%� U�ٗ��f�W
���`�w,e�ٔZϫ���^�u��j�"���8�@<p;���"�Q�%!T��Lv��
9�D����T�6S�Q�F��4�퐵���G �e����)�/�ǽ#�j��j(��S����:�T}����el�V���d)|���^K.��Ұ�Z��CP�-�	�������&��OXa ���@�X�HAo�>��#�C��g1��8V�Lv��u/�گE!Vg�gx�V,��X}��H�x:���^@�x#K��P���>�K��g�G�1�F]E�N���غ��J-T
��R*Ƥ����ޑ��Z���j��8�?���j����񩸰�;$�D[���*�q?-GB{ٙ���o���B��=O��zM��*��3�i�����Be/�*U0��dt9����L�WH���R�����76usHJ��I����İ,D�G�>qG��]��`�c|&��"��9�S~�ڍ�������@��ܟ_c䶸w	�9���r�i��j�qA�!���#���N��b�A(�jD�0�TNËzi�X�o����Z������/0؉(��{ש��D�ٓ ��Ð����N�H�� �;�,�������tf���R�ɐ/��u�9��8����[&�Zii�ץ�
�����]��8=l���4x\�w�J�O���"{M�`�`�OLߴDB�P2�� 2^t�������YMF)�P!�T�:}�U�m
O��\�o����
U2# Q�-�H{�0I>��\���Y?Yo�������mBRx~	�*^�X!x�42-u'��'c��=Z:�nĂ�W�<h�������ti!�	�]��H��\��_�nA��y�Ɨ�t���i�YX�«c����	����'F����C�hz^[���EP,����<qxN�h��/������/M����m �tb��	_�aIk�REk�=VJ�Gfzs�U��o��=�4��2Yn�܆d1��-\"	�Ł�r�n9D���O�T7[ ��y.
 ��sJ��ǛM]�/�".9�#�1�Oӛ�m�p�����tb �:U��\�H�I��4Y?�T��#����(�l�Xgk�:2⟰(����SNWM�6��~���o�dr>�YU)J3�C]vZq��9�|�(҉Ѕ�l������$^�n�L��w`�����&]�[��C���a����H���k^���c2)��B5#�<���@
�u�+v7�����ͿV���J�A=/���kI��kc5�x�c%C��뿘�y�z��d*�C�:~�K���	���kl������<������j��9j<����Pk�}�6��
k���R�ӵ=�&�wd<��#�b��-s;���c��*���� �������/[��pJ!ir"��* �"�/B���sv"n��0�
�[zG�3��e�F�+�κ�.(e�2�q)�tU���ҕ��c�Y�~�)�))��MҲf�Xh��yS	���v뇨�����g��"����u�GK6Yw.�A�Wjj}����+�C��܇|�H'��w/��l��%� W.��s� Q�o@���vT������8��}Bt�.�KHi(%v
V��K�r:��Iْ�]��;��������Rs5=�e^C��o�����f�����T�6���@��ud�<��u� A�V&D�؃�P���J׶滁5g���Z޾�Uz���Σ�S}�5)��d���ZRc��!zoE�A+b��rU+- 8�z�t��"���\�0L/Z%��
�)�����(,�E�U|�,��0��GЦ.��;��U*=0�q��?Q�4x}�J�6�J[�r��Z��a���ԺmǉNd#&	�������I�	�
���	�wD]S�_H�7��tNA�\���nFj��W3�g�[�B���?nO;^P�A	"��b&R�uBPq��n�����T�ԡ��C�q�x�Q���<M��A,�;F.��i�1s(��!B��G�S����q���6�	g�p�'#���Kdsn6��⚁e(T�l��鉥��d�k~�<D 꽿zF������-��>�;�t<��zn+w0�"�
�����3��.�PF/|>���e�  R��s�p���p?�!�,eS��;��ѰC�X�!$��f�e��/C`�r�����9]#�y��R.}a�ϝH�T�8�a���-����f���ݙ�m6��W�"��/���v��l�|�x�b3�z�刈/P�|ԩ�~(
jKe�.�ͳI��r(w�л��厖	J@z�*Xu:W�����V��?�Ȗ �kh87�X3�\����%����B��*J�&�k�U����Ϳ���QUT{�",�;��N�'",��O
���y�v��ߧ{����a	�wi���#:]����b�G-[���e�3�|=J�'~�R�˺v�Ò�-l�cP��M�9�D��$|���.��B��oԵЈ��P�)f��U���/���>��h}}e��V�KZ|�fʏ@�0�i��}��/��.J^@�L>�o �2��9d)#-
���1��U����-��� �ឿ�5��P���e�u}B<7`b�ܜ�ˮ9�*��M��}��Mc��"��t+�B���s�iRO�S~b5�^�KfZX��f�=j�6��.,�z�+
��WonՈ���z.� ø�lX,Bv^�nÌ�i�g{q��LJ�=u��z|`�3�n�̿#�;�-^O���_��˥�$���eU��o-W�y���*��a�x�,ϳP��'�B1�p�S.k�WJ�&o^=W�J�
^v{��(ud�-����.d�&��N4H6Af�8@��p����U����^+h���,f7�:�6���Xw�E��������:f�D`\�����t�/�	��I��Z�'|��1{���A6v�g��1~=��=�L����}�[}!�R���Q"��Kb!TEd1ZD���`�C%g��O[�Z��e'�G֍�}G��qh���3+�}L^4~('�ZWy�y��� S�1!J�-D%�a�7��b���@Ai%�.ph�cv9�!@�U�P�2~���8P ��;c`��CPٹU�=�"T:�_�̈�#��yz�e7�G*��4�W��;�_7*��7qY�fr���ǽ����6�aD���(/�-���'���q�?D_q/�l�x]����:��llĄ���zs�J0�2u%/�>�mck�#����f����o�Q�3��萅v2�y��D�Gc�>��Y��$�c���ٴ����_U-C,�񅟃�H��a��P���:��>����rq���"�i5�ǹ�'�D�E2��'�L�ꅔ�+�ȥJ:�І�^71��η(8�G�1�~���l'�-O �8�k%�c�}6��,����8�g[��SKAP�	4�����q����r}�Y����uc򰦺��<�\K�,[�L�T1�^��g�3R���Ü�`��CR7�Z)�&�TdYA�Q�������.�,���

�9������3¬ (v�i��Z��9e �3;Q����Q��p�������a��
����=8�A�Zǰ~+=�7���GW���DP*��i㮠I�V(hc1��:83\��f����A���y~�~Q��ʐ�-������l�(�t~h+�-���[k�}=E��d��� �9����hpl��'�F �~�7�j�8([���z}�]
��u�UU����}jN%+!����f7�IƦ�%DN���B�D�v����֩�A54�N���L�#	�ʴR��L��5�Y���«�2:�22ey�B���S�J�F�E�F�(��<����ǈ�`���6�q,a7,���=��u�D���N��$����?���\豝��E*���#��jR�}�WI���Gux���L�R{��%���tN�)z��4"?������p�E�c�y��DL�8��	���J�`I*^��=�i�hfN=M�y�z���z�b�k}9�w�;2 �����NS1�aZZmK���[�8ㅁ�1�E���G�����f8����P,�	櫏/S���<�`sg
cN4(K3.�Zf8-'���W��Ku�0�=�Hb��Ï�y�ɯ���J�,�.��0gZM�%����D��+%��T�2���h���F�řuV�/��'ܬ.��[��Vyxe�s'��l'K�[k_�ӭ#?�,� �f�U��3\�DTJ�Dt�'�xZ�*+��	���D�+ZT<רj�)+��$�Ȝ3�_f�5,���Y؞��s���)$V��uU��J�z�E�d�~�}ĳ#��N�ۨ1tSF�`�� ��\�c��~�1S���x���#9�{�!���72U�w�<�pj����Z�>��8��l6D�������L�'K�q���VA-ܯ��Âux�B�$<%�Wv"�`�S6˼��ޙ�����Ϙp5 �f1n�$J��f�̱������6@v|x! T3f�4���IC@������.p��4�p��4�<r�H�(��p���!�"����zޖ�
�2����$��؄�ʎX(V��Y4s`�@J��RS��{U���~I��=lX����͇
����Q��7�������7�p
^�:�ME�"�N�n)��:�Qҷ���n�e���J�ђ�Ҏ�<tN����i.0�]���Q��z�ݮ ����pd�rT��$� �ڮg|�r�N��@,���{�������3�?E�-(tH&$�� q]q|s��B�+-���p'u�G�C�sn���x��d.�N���(y��R�>h^9۟*D-q�x�{&*J�����x���cS2���B)��|ۚ���L+�(m�k]�/T(+=�V�i ��� �kZ(?��Q7�Ԣ������_p�4g�|��$�G0����<.��J�/[�
��<0��؄hGG᭙�+���c���	f[@ߔf3����Ǻl:��k8�{�M��0�8|���]fO�9!�-F!#�w7��X���]��O����5��ң(�G��2�~���I�_6��	��R�����1?� ��	��W�i��~d�����a�In�U�\�|��_e� ���7���&��79D�ۺ�2n�;�<ׯ�a�C�UdV`������1됩��Q9>�ar��(O;+�"/�L��ƚ ����NhvN�6>���4'���-�����4&G�us�!7��
h�R;�2}W��G��<����3��:�fM̔�o(�3hd=#H������bϝ#n~�Ф���1Y����@>��Z~�e���v�����	 �R��`��%C�5|6���*>оd�z%k�1�y{��:��nwϟ�#����3��?n>�r\�]�U�I��E{4�c��଴G��2�7o�T��'�< ���j.I����z��1�R�Ӏ��.�_���t�zΐ�2��ž��5����@��iS&��!����F�~�ƆF5f�sOi���8��_����ĖTt�9��Ʉ�����ǋ�-�m�sl�)|��i*d\N�,�z 3n�-�N��%ӦBNt_�h��N{ ���i	F��[�,Oz�5�7R�, �+�aLŻ����{A��K#�����n�+ǎ��,4��+d?,;��=F}
�����e��Nip�
?�Ω��]���e��>�& �h�D�"κn��y)z���H�Br�/���ӭ���~e�Y�3ϊ�������G٧�\�p��M�lP"����S̓�\�(h�B��`�~�\�r�]R����,8�������TZS�@!kэ�]�J��gG��YW	"E���"Ɏ�iն�ZQR8J|q���>��jF$*�h�#��!�%p�aٍ�)/�>Ne;]�ٰx�?U���"L��iUj7u��GXd��WA;��$"�"X+2��ի��ux�S�[�OE���'K���ݣ���b6���p�*W����X
�?�M�2O��M�E%F�:YF:��pxf�����u�׃�!UQ\�Ѩ�v���i1�\dH1� V�����y)3}��v[+tfI�+�vΝ������l�V�񓍕 x��N �#i����@|]#�٘_�z��W�&��Um)[����Nӎ���qd�pغ���ee(�Drqo	�1Z��쥸���v�E5?���7>=�ՠ ���Z�~R�*�橌�r�Y�i���r{��$_��q��w���W��QTX����5���ED�?/;����z��~� d(T���C4M�X�+��}�B��.N�U�8��B"�?�Ҏ�D��R`"t���+\E1�������(� ��;:��|�χ�c�Q�u����Q���Ӄ�9[��o��e�8�P�	���bJ��uAl�����b�4�t�ߐk�y�Kb2o��m��VB�9�m�`�9Ё�,����j�ة;�<��NT;�%�]��4�ď0�e����*u�4&犎�j�@��ۜ�;�wk�:��qO���q���	��_�K� O��o ����R\<�+�Cn}������&�+�n�̓Q��n2$��p�Y��`������h���X���G�J��+;�&}��'�d��%��^���F�H
�J�8W:��Z�˾�iÒ�.�Ap%��s��9��P�G�׌���F��$P�jRR_��]��Q;E�t���89��7uE��/�<DDc�ď�K�o� ��	��K�[H�u�TA}h��m?�{7�'�
��;�er~�Ōވ�?�	y�䃞,�_�y��[g�oS%��ɷ��a�jk݆]�q	���TT>o��z�{4(���N ���X�K�d�ӊ�,Â�k�㋭�j������,��0��'-�ج��B�X�ϐ�(����,�m��}d�V�'N t�*ݙ��O�':c1i<�0ލ-���K�t��B".�b�_F2�8��_C^M���{`z�'#G=s���zH��A���������$���� ���I���]��e�*�}O�倀����Nx�.@8����w�Q��t���A���e<��1�M����Z��akKD�m��� P#ןʌ��{`T�t��yW �!�(,^n��q����@D��q݁��P/�A_p��^��}B���uP�� ����/Y)�����2
l��'XJn�6�����=
!ƒ�f����G1�F�I���Hr�p�&Q��I�g�g�񡏒��%��4�7AY�ikNdĹe����$�f�&���-�!��=B~�u'[��S��w�g�@GU�Ee_�?5�[��	�]�nݏ_V��8���JPC��;�\�je��5��D+{h�k���<��\�	?�[н &@�j\����3,����	y�����ִ��/w[�!�3�0�0Y�4 :�DQ�Y���C�/$|�>L������M?]:0�w}l0%�r�%l1Pw�k[������zZ� �P�Yc^��}|�)P�@�'��y	X�|��V̙�xN�C�3W�^:��d=�QW%,�WJ�d�SY�G��VOW�ٰc���P 0�^�0U�ޱ�Ԣ���A��guꑞx.��U�c�>f8�6�����jbH�wXQ��\�i�S����\o5�����A�9�)�\�lPj��BL��ϔ�U'�'�}�^���S�a�_c*ݙ��3�:@����$�$\kUF��=:w��u���P�6�c��Yt:k�9�`���/��p��m�S���� ��*�PH�	�b4�:��D�3~�Tu����le�������f�D��G�1�|���U�9��W��l؅|; �?����Rk���wܔ���wt�Ne��S
��-�ڡV#M�#�yyp�ē�Sa|�FK�Q�N��s�v�-��ւ8���N�C7q����c�j�+.6#E?��d7��*L��/�݋%�ܛ\nH��|SA%:��W���T�C�[n5��E���!ѐ�Lq�g ~Fc�
�h�̦i�<1r(��˞V��Ȳ��S�z�^�����4�d⎂@��&~��EJ��K�m�t��V���X]ݡޛ>�A:!�^kg>@,�N%�{��	4�<��xS���>�g��d�s�p��ț<�ʲ�݀s\^�P�x>h�j�cj3��c�k7 �OR���/Y�FW�N0��[��D��~o�U&h�h�3j���&���@�աӣЇH���a��Q7���\V�t�#g^ ��sgQ�.�F}z Ol�4��-$h�[��T�V�o���oӣ����_�5 �LʂGi"���6gS��p�jkAf��X���	��&�|�=��:8��� E��47��s1�}L�h�iP8#f�X�q`���">���=�*��E�'�:��Q{�xv�0�E�+"]��F�Qu@�_h�bt%�dJ�,��M�r�˺ؐ6�&%��QS>��vTt���h@�B����Ĭs��eB��N!`x�p�'?|��Þ�£c%��y�l�OV�Ά {X�Mb���Kj(�*�dv���4����+����|�4�#��g�Q"�63���Mpp	j+D3����۰� a*:����B3��F���`d�E]���jt�DKK�f�ӯ_�UܞS�$�-ʟ�_�c
C��@;��s$c���n���W���o0X�6��,.)��?��^*�����D߼|���ɖ����5֐\W��~��������m�4%�k(&"�X'@��3�|�Tv���Dn=q(�A���+�ba���J�#g���Xb��v�
h(&�2�<�h���ȸR�+�^��ikj3邙 0b��д*�E��36����zҗf�M6�$����� �$���}}�*���^@����îЁW�O���4�;���\T�%�]��x�.�F�V��Iի��Kz���ԫ�Կ����h�[���E��S�ٞ�<�A��$�BF�DC�@_
)��M#�S`�����=���lרV�YC�H���5�r�M��ʍvs���vٞ��8%m�,�����)���⛚�D"g�%i�c`����o�T �U,�'��j��[�x�4�s�|��S�J�{u��	h��p��������G߄R�Ì_$-)'9�\�5���g�;���׺�«�C)�[��̸�ߠH�2��zf�y��@U��?G�g
�cubF����QY9�<x�BsX�>����Q\�-lm(�]��[�8
�8�R���v�j��w�pCw+�b4<��%n+mSQ�U�Iu�ځ�gC�<=�NV99�bZ#�9��9%%��Wq����JB�B�:5� �}�D�1���b+̨��g×@�@H[���c�8��_m���74�+��~�yK���۹>�5���R�L���O�m<�C���t?��: |�t�|�U+���K)m���P�c��
��8J�+ioW߆	7�
(�:��yb(�\�{nP�S���
Q��5��e�����|\�r�h�@��8���96���[�zG���U&�b�O<�8��,v���
 ��g��S��o�5Ad<ظ�ro�U���倒>�ϗr��%��S�l*�-ʓ}A$P��[�(���e�Z�S��˓ݾ����ʵ�[ۼ8z���7h�����6�{��_�T&	v��x���Ö;�2�&QW9���Ŝ* ����}Ѐ4�at��V�	l�:@Y���P����c-��-	�{S��"��_䚿��j��<!�&���2
"2�����PVC�h~ Ű:�D����C��D`��fy��������;�鴅*�h*��tEF��[��@����7�0���y�j����J��2�pU�/��]dm�� �~�v�	f����I���
��Q�?�3��?8W���rY�᠘���fc����	�=��F���֘bO��o�"<9��~�����)A�sߏ�Z��}<��Vly
�4.� B���H��ЃԺ0�?8�WC?R��;�ku��2�Sl��bh��r����(�'au�p��*�1�
�M��k�;��_�O�bMe~~��>����+�Ƀ���|M�$��z,'��ap��DD�0GM���6�-��
�Z��@^MQ��B
�8��L(��Ȗ}�o�5���D/�� �v��9�E3r�aC��p1��	p�-�]����#�:�Z�����:���]n	�}w� �����8�)��6V�WR�_�!j��;�EL�6�?K�b��$�A��~+O�=��9x�m�j�v�V��3)G^�oGj�T�:-�M-�uTW����!�#X!θ�+Fv'IJ��(���ba�?0�Q]����=g���+��&������_Y؏:���<4��
tMW�Y�_E�ė���o�7�aI1VM������(�L�!��r�IʂN����a?~�.|�C$ѩ�.,�p�q������$�'�&���UӬ����%2wcqҎT�,�B��?l�J�q�B� �'w������� 9k�Z$����b2�.s�ٴ I�T�����@�6�~Z���\AW�bQ4K77fc��.s؀{������ə��-~̗��7��z��,j�gQ�3�v�]�?
z�c(i�����7��F��@cߴ�4�5�d���ĉM2.d��z_�ľ�l�L!U��6�A�ݜg����@TeK��uF�i,�R���T�z���W��<W0րp����q�Le�T��,"�WS1�
z���߹f`[�e�m�d����y�<F�8d�ݹ���+�g	�kk�2��f�I�j�ð�]�0��#�I�Ă�������(��F?v�-�j�8[y]����U#� M(b.W�u��GlKZP\b��d�P��]Ge��Kn��bRGI���8�zƬ�A�+`Q�#������^�(���\ji��P�I�6D�>ЎC�TB/���
�hZ�x��hڹ;9�%�9�lxޟ��c?toF(�6�Kq���\�?�X� �M�ئ��X`@*Z� ��@
�|�'��0�sՐ��PBS���6��2�RfӢ�!�P�$1!G�����Z�$�߶�^��||y���)T�\��c���P�H7�4|�ә�$Ϩ�Y��t��7�[U���ː�-�̾�x1��i���@�`��QZh������5���Uz}4��[̕	�������=I������'U�{�/*��U��b�F���Kh��]�lѕ>���Q ��F%)�wId;М��/��h3[2F�$���E����al�>L��s[f������E&HZ���d�/x�"��ޞУPtb�����4�U�Zaj�g �]�ٝ�fz���H."�hbL>/�u�Q�J{?g�AG���F���wv���<�9���FeI��
���d�c�`i���l�r���G�$�#���n��F��W�Eo]��^�\��#k�H�ӐS���='�?U��)��VX-�@�6���λ�B*}+Q��T��9�kQ��w��o�&������8X
j�?�]�߷�����b�9d�:$m���vdPp�|�ؼ ��d����oR�[U��O�r�S6l[
��c�`�����hߤYL�����i�*4�Th����4���H�.
M~�x�KJ���~0K���G���:��
�&�Y���2����hע��»tEvȏ~�$9��~�-g����p����`宥���G��㎲;1��URw-1�C�����/i7��S�dC>����Es��/G>�|�/��AyLA�i\���W�����y�^^��"�6�&��
E�U���[3�NA�Ǽ�t0����)R������]�����7�q��R�����:]�X�x�E�u�'IF�|�/7��z0�)���)��e�eYb��.El!�d�i�S��������[���z8�U���0G:}������w�@�1�#X�W'_x�X]�;��{����|]�y�[���z�{�^y)�4倆���Y���45���{��]t�Ak9�H�$y�KE�ۥ����x��K��t�-��2Yo;Hw�p�U��ep�y�JA��C5@��Q�#1�!�����ԝ�&lWn�Y��<)P�=�~��-ӆ�9��"�Y��VbF��.2����o�\I��������׬sr�+G��`��Zg�:��4$�ٌ&��̍	ÕQ(QA��Ԓ���ݢ�/(�U�� �O�PNA���Xk�!/�uAhc#A��tMz5~��9g���#��Zִ�f�ƈ]�à1A۽��*A��c��+Q7�,�Z/����� �&�Xk�֯J^�|֌�9�%C��}��])r����G�'~w�z�C�h;e�&��v�u���?��F����9���<Ŭcd{G�=��Sh�c�}_�Q]B��� dN�Ċ$y$�Z�d^�j��� VS�J'��3$ʝ2�z$��]�h���89��{�^���,c�=Ȋ��x����m�L���	���;pCOD.�ƾ1��:�e�������uɱ�T��������s5���Y�?����dY�9������A��hT�u8��/	΋A�־ǮO�������w����XfFAP��r�]��u9+�P^��$��z��o�n�=ג��Z�0�U�ч����(�%0��wA��xm�7����LR��X�چe�y7Q�"�\%�;�������g�Ŷ���P�%�ӵ��?8��[���P�������Si^�`����@=QYT6��Eʏs��9~h����v�Ȁ��!�b(�}�㍞��/�8��j�F��}�5P���e�d�%�J@�o��N>.��Bw8���Д:(%U���2~I�F��	P1݋���b�H�/KW�?P��Z)B鏨�.�;HDaߐ���ddU�����~nh��#�:�B�9�0i�|�/���yq�$ǝ�1ҏ��]�\��)	 ��_Q���`D�����|ct	o�Ϲ��D^��~�r��SU�y w����G�	��S�����=���4���Rws�_��Z�Șx˖���
�\3�^e�m���=��_��ĉ'Q	c�௶���U�F#�rEl�V�,4)����B�e!#�����RK�t�v5c��2H=���Μ!)�ߢ�h*�&�+��H����X%룏>�YϹk��B譯��o�k1ȵ��CՊg��|�������F�����qD��ٴxY��絒�`��:�c�G#��t�&�%�D�-m�'sd2$�B�a�;���w�`�}A0>� �p�U��CԷ����[�N�{/�4u#�J��W�\�\�>%7�9�)��]��S'*���Uk��ޟ2�E%�9w8��XM�̒2v1�+z��n�e!ɓh�h��,-�Z�,��.p�w�cp�v?y.�@tC3 G���M�]�2����r�UMҧ��*�����8Q��:��p�AQ�ϝv��X�sb���>0]��֪oޔ����)�?��YÇ��+ؗs�F�:�Aʰ�Q��u<�,���u��w E�&C�����q��kb �`����X���~M�˅up���%��v9�I�R���	\;6�s�}�2m�('?��}L`jR+�
8zC� � �)�x�þA:�C�+.��"�v���9Bz��{���t��`����Mz�Z��ڰ��,��P�I:������j�(X�Zԧ6��g���5,K�JN�8�m"��g�_�b���*,��N���3�J�?���7��_���xt�F�a��f��͝͆ ���ZT��>q&�>���g�9�õ���WV}�Ѭr���%1&��6���Q�m�a�y&L(����	��,e��S���Woi�{J��&MhPUu���8"4���'Zx����]������W^�z�44�x tL�uݳޞ��#�/;��:��r`��v��	�� ���)V��`���o�����8��;d�Ƭ��)�Ɖ���� �N���P�.7r�9�6N����Ks;��]��,%�I�ˬ]�<.������:+��@�(s[>�b��uC�ruk�<(Iњ����q��gs��vij�+fW))�9�߬�LM�^��|��g"�?���JkI���E���b�{�~� �9Qᅋu3��y/k�8�����<��~T�z� �� s#Y��{�51�f����>��U�? >�頴O�:�4@�C�v��0��ٓR�4F�JKb�,Z/b��`S���A����l��x:U&�,zF4����}�8��OX~�Ê�������1$�r��T�R�V5��?>,l�-�/� #��z�N]E{T�R�M˚��C-��
D����^������B���(��C�~b��Ω����g���:�ois��+~D&y��i���֡]gg2`�О�?3����	t�e���_u�3�lV�d�E��o��B�{��^+��v�X��ty�7�J�TK�Xм�g�m�/W��vر�dz�_G����;ρgW�g��^	� #^��)�A�ةx�Dw���8;��>7����^��sHvJsQN�:�@	�3�s�jʷ�	g�l��&�����D�Y��%�E���s���ٓ'�h�����V�5=�,5�gh�%Ӏ2�33��y�	�}c�C��XI�$5F�hx���TYܞ�����>>���^�=��jǮ�bsg}����GU�l������<~n�~6�B��-��Κp����d�_#0�G(K�u�o~�8el�iOY}n�SM�U��rbs�����B�N�3��]�������9�@֤�X�[W�x(̠�8):U��jZ�mրy:���
���A#ѻv��T�W܏�7"�:'20�:GQ�u��G����ʀb����7QҰ$Q��g�"�TI�!:ZH�Q���Z��@�v'f��|1ß���$`�����b�ӎ�,�&m�>%�����,�;M�__��e�Hi�[�6B��Rx#������+��J���NŖ���?�_�e4�"���뷻���
`,����3_ҡ��7��fIi�|�λ�C��"�>�*�BZ,Ibl�X���E��,���W�h��JM�o�mn%��ʬ�����`Y��HI���7��m�rO�g}w��N1�|�@�{t�U��!���&��b��Ǩ��R;Zɇ#vG$���Jg�͋�S+������
P�=��ł�h!�?��"�5���*s�Y'�w�:4c���)������Z�o&ϼ}ކ�譳UAn���;c��$�P&Vfk������2m��aY�jT�#����!)bV��������˔��Tp�-����:�&5;NQx��H�!���^�ҏ�ϼ�ADNRO�N�1��wZ-1� �\0�t�4>�.Iߊ���w�ݺ�[���a�ʝv�F�m�k���6��y�m����T���l�R��D㶆Γf�m��q�}:��Y��U�� �T����V�9��{Ig"��w��˳�_[�hb�#��x]ؿ-�`�j��6/	�&�<����5��0ige5m�O%���|��#�/� �آڈ�޹IW�,חU���� ��*t�YT rx��R��A
�㫠�ݢ�`U²����eC&y^`�<�;����*�o��f�ߧЮ�	�?�)a
S�L�h�61v���^%�d=���]t�H:�Zt5x/��a��U����N�u����fbT���]H.J-�^��0�,�>��<8�w�d$����:*�Z_�u|�XC�~Г�וK�ͰV{C�!�j�'�}W������ŏ��H�/���� 23�U˯imޮQ?��x65I�.2�Y� �s�.�d��&�%�}���E�&��U�+�TgR���\h@撨�Oi$�q�j�>�ps7bI�)�F�'"|Q.\tbt�{�m3x����TT�LϪV�^��D�:$a����>,��Y[�zR�%��FA�2T���{b��(���{����|�⽲�[u��H5Y���m���HR�g{@9��U�;��DvE�L���~�~��e��@��4���,��3\Be���(�^�����i��P�+�?�����_"��th�G�_��~N��+��ڸy
B{S��?�ʤ�ԙl~A�����漳\Q��RBuq�-�h�t(g1b5F�m�^�H�r���g-���Si0�ӕ�CA��.�h���!"\Ŀp30�~&C�¯�s!�r����Ux���}��l~3���q�~�D���]M�m�`��>�r��%w�.I��T�_�ap ��HqAl���^}���k���*^�Î�J�Żo������z�w4��:��X��E�'���h�'���c#��eH�?Ǳ�RMk͔�F��7�gB#g97;�>�9�o)�����Qm��^��dǿ��i�L/(��^ �*��F�@���;+Ϙ��5O��G�]�yn�e�lv�I�1N�	(q6q����lDa��NT�vE��u��yfڞ�B�g-�� kG%����;Y`���NU�zڔ]��C���'��6]d�Y�<�|u����_�eqEY�:-�pL#�5�^y�KJ��
���h�w+`e@{ɗ�����g����3����tB���*��a��LW���(�ֆ2��	-5���>a�6<u�k���o�q�G��1�DW|(V��
���@VɌ���.������!�E��L���U]nIJ����w�S�V��Z�n� m��i�z	4��v�n�e�ʝ���i��X�J�9�+E�e�Z2{HLѺ#X�w/�v��Z�MJu�����\�0u���;��2��*~�R<Ã������V���~�_�r�ʫ��<"W�Ⱥő�F=i���<��A�{�{Xp��8�c��#�� c��MY�=�%����X� �+�9w��сy[K����};�d���cz�;�E+.w�l$]�{�WU��W�5x����D#^-�B��riك�����bajE�~�r�yK<�Α

�5����=(/ԷҶ��6h�[ ����僶Yɽ��Ӄ>=������(�~���_�O��I�@�D��X'arD��d߫�5~�ߔ%>��Z�����4��`ؘ:Bl�p[��flbg�;&���:`�!W�	�5Ձ2t�O���HH�AP�ōi�D��MHGVU|'������4�Qů�U�}L�=�M4k���`��7e4^�A�ߦB�b[�(���V;|���
f��[���S�/,��gΘT���\�E<Go���qI�>�O͚��[s������4^YFjކ�ȅj�".�v��L_<NF���F/?p�:�b��%�=R��H�|d�lW��.��K箺-jFq�����L)%�b���祮p#�<�>�{�%�H�ꩬ�,�^.a��D�>�!��#.��Ԝvp�3 A�<C4��!;�*�N���(��B�W�a:����Ŧ�|Z���O�F��;_�<���`��[B`�����/�� g��T܎����!D/�1]����M�󉷛j�V�˖��e����}5y�$%��l��P�&,�Y,���!�/�'�Q����Z$ǹ|UXz�� dЪ=��M˘߄���ļ��3{�=���!|횧���Dq��\�~�t���a��{8��������R�N��-ˎ䩇�"d��L 5g}��"F�lG-U�fd!�������#vh�O~S]Zw�;�eJe���6��9�>4�<��Q@�?b!5�&���6���"��t�^�H�����3��m��Ȧ�J��d"���ֱv(+����M3�f��+�VN������I�s�&�\K�SE�Y�S���Y�;L{�����z��� �=ϩ��Dt҉b��Y��q��n��VazP;����L�/"�4�\=����q��.=d�� ���.�{�Cj����8f/��0Z�0���ӹ��1H���E�b����!�UL���[mҔ�i�+G�p�=��d=y R�֬;�W�E3xa%��吉�F���@�a,�I����x($��&�os!�)z�B�:�Mi�"0��}��G���?L=0<��`N{B0q���lnl�����1��Ԍ�V���(I���{6�����^�V��j5���@�0������g&	�4~$��@��7D�d�&}���O+Q4�O�g���g%2la<����z��m��S8԰��X�ԭжt�;S�&�[.W�m!��%T�ܗ'��
��z�CZ#
v�I�����~ی�G����y�bm���$���>6�Ch�ғ^ ��l���WE���!Q�E��"? Cǥ�↵ɺ�$$N��Q�����^�gG���U���e�1�">:�Ȇ
���@r��b�X��������F��y&�m
J��#v1WHêw�rT��"~�����uc���C�ҫE�Tҫ^AW��0�kIY������ �+��;r��?e�����D*p���7mzD��N�cAǉ��u��_�j��'��l�S0Q��̬3��x�F�^nfˆ3�Fa�d�f:F��V�@e�cN�~���"b*T%T�@�gF�[�:n�|ı~X���x�!fD)�q������̰b���8�Sg��Q��$3rl=% �]aA;����U	��~ԠJ����^%��F�[����#��m�P�6
��e�:T��м�c垤,�Mq�#6'�k���Q��������1�\�)VY��z͘*���*�8�?���Q|�jX���K�9J���޺7��ķ��:*K���gn	��E��)6\y�����կ����LU�q��Ӂ���I
�B�q�S|�2�I�\���"�� iҟYZmn�EH�,�4=m�y�iO�� ���j3k��C������IOW�6�2΀��4�_P�z��)v�;+K/���(���9����m�c��ȏ��2Zr�y�ǔ`���5[L��X�)\� ��8�Dt�?l�;-�)�p׹I�ul�G�n`e�fzl8��M\먍���ᘛ:d9�d��������П;Կ���R����L���Ui�O��m �9[x6�GOPy1=T�	G��G��:Ş5!�"J��d�W�f��w3�wv
�ΎN/\ۋ�'��3��W�c���@���Vtvh�� �%��x�,�,�D�7IOΘ�.�����1ӵ��ʣ���&��x�n�~RI'tkJ�����zֈ���6��lg2�2�6������~��+q�H�6���}�.8(�ɘ��R�����a`*�:gj�����fL?�Bɮ�-�<+�(0�?�C����=�7֐�z�_�!p ��à���a@�?���H�n�yI����'��+������pxqL_�p���G�iS����a-L��Ș����aD���ֶ�2��?|E�5����P��Spr+����>.Zޔn��v!Җp#��m��޸���Vq[��a���ME��q�O,�����}�١��	���窗j����xWG��W�s�J��t?�!���	K@C�ꥠ�����R걈�|�)P���p��5��XD_p,`�K�SB{Z����)�i�}���WaE��|�����,��3=q�z���'��zpD�N1��xeQCT�XF�X�%�Ȝ�yP���r��a&B��0�髹�9~��j�^�2�2c��9Hwħ�Qp����EQ���HlV���جsg5D�:0耎z��EOmR;�lX��d��6��T�S���QZ;��E�Q��nc�̲%D���.��)��]�w�gZ����2Eg�B���vu��cQ?
��'=�\�:�z��8�Vl;���_ͻw=�ј�J��镊�uO�8���V01;� ���	Y�w��~�ԼQa�7{.���}���~Zz�IG���S
x�����R���`)�t3��Y]�*y~�{�R/����j-~��Q�xsu&��.� ����,����dЋi������)��ޱ�6qD�Q�.4\�בi��rq;��W�e��U����s��_E�C��a'�6B/�]�6�	�VǶQ��=�ɐ����J.�o;��i�^�}����'p��U#�ut�
 lSD�l�j����CR��b��������<k\H{:�Q��Ǔ%���o{��I ����h
aPA���#o����|?.�PeO��7x��ӃGf�D������N�uθC
���
��b#�(���_?�OP�%�G5)�	�^�/��(�w�ʲ�` ѵ��(���K�>,� X����֒�X A[4�<�w��Dd�����_��D�2+3�֟5�b����ǉI�v��!��<��?�s��H2Y�!�C��Ly��u�L�D��ѥRmm]'O\�=�L��Λ��1	�Ȯ���y��������{�������˶!�wm���&@>�2.���2��I �[����c0z4�~6�����sQ�(,/"c:����M�ZH�
M���g�YS���P��\
a���W�(��A~�b���^z�"��1������Bk�J����xg��@�>ԅ4c����mi?�Ń�R�{xUH�u�\!��|��T���0npL2������0�Ġ�SΗ*�o�� ����)a��ӂ�zI�����x��ҏ���i���1;r-��@������|�RJ��O��c���ahK��6���@N�|�į���]	IR��AP�<N������S���X7���b�>��ˎB���x�j������ �D �5%on��)ST��s$�ą�!f�|H$3J���x�ͬ�}���"��kn����'`T1w��\9�7�C����_}�&��2U�� ��>g!�!���z>�X�
���w��\@��B��Q����
x�?�=�`���uyŴ���S
�
|�RX��^%�G�(}�*�m��B/_�s�wv
|���Y�7l�H����	\���#�#,���e�%��
�_�P�;d�"���I�^]��r�,��@�Ko?��0�g��; �v��C<39FY
�k7��ɑ���}=���t��k�%�ڜ����l����?g���ޤ����S̭A~�
�a9Yɞ��oW$O���0z�f�7չ�)t9��1��	�N:��JW�3��m��{(j�H�p��|�L�@�9������sH���(�i�K���/�^�Iǽ0E���	r�M�s�6�5�w�,�r[@�O��4�C�ee��"��B���L���er�,ϓN|l��椚8�š���qQ4(��m����l���h33��Š0ݥ�%�3z�[)�9f��i��CE��0.���;�9-���/C��@J�k�whVB�q�cv�o���Fp�О5�z��q�O7RH~qA��h�g�:�l�"�U�}m?j�1�Ki���K�e[� ��������-7ޯA���Qy�;0�ZJ�� ��]V��kC����¾�(�qy|�+�~9�wv��J��=���à�mG7��F�\ 4��_e�*����.�\r�Y<��	�H� D�Ll �����Z{'�nb��<y���Nx���_V�Cvnԉ�Npp��`��]�.#��yO `�����t �0'&S��Ko�Y��HGQě�&u���1��,?5���/�Gk��U	�RǦN�F�/��話6;�;,N�,��p���\+���m�+�.��p�_�'�8��O�\� ����0k��q����������VfJ�60Q=�.!����,�j�f�������'�{�@��.�N�ڮTq�<w�Wr������y$�o��S�RV��>H�cB"t� �<�������#������߹�xd���a�! 0���땅fv�S鬱?,��*�yn.�F�L�J�D|9�B�}.M�H�ig�2q'ڼ� �j������&��Q
U��C�I����C�v�u�g��7���|o���hlU�`�	�{�X�zl>��yGOx�P@�S�I�h[����b����f�Ch��o��#��t������sxdpҒz�q}t�L��}_訮�z�!SKk9���,����� };���[��)&Z5�s�Pk�km=(O{e�����WF�x�me�1O�LL��bJ��
�KPuB\\%/���f}SA�-=g�q	!d�\5B'�9})����]9�s����{E��~P�1���*l��+�ψ���Y����iL|A�{�3�ڬ��x�Rg4[�b���)�vE.����"���ۨz�����}Ⱪ{�(�Z[�$�Ѫ⻺��4h���;F�bHQp|�Y�K���6��c�J�l���`�bH;�i�c}a�ө��.�77���x�F��b��Jx&�*�(��x�M�>�<�Q����\;� ��+���R$���yidA�4$�ԍ�p�SO�M�%�ir٥i�����
s4
fxZ�+�
�J3G�L�ؕ@�o��j֟��W��30�5��Ay�쨪�Oh�, ���ݾ����;0�σ*�p�f6��-Ī�ح>[���N[�Z�g\d�9CO�+�9a�I.A���Sb[�1Š�����������G}�عJL����a�^���bݚ��(������{�<.W�9�t�&��A�~�r6�|�,����~����^��g(��$i��,��k�~������|�~;r�֭)	N)ޖ۶s�sTs4N���c�ϐ�k�ga��WIs>+��SR��Cf�p2�a��"G&r�����U���kWӄ����*r��ͺ�S��b��5LKa�_7�|䈠��
���\��O�	�_@$Q����ӟ�N���Ы�1�k��B*��_��RE�2�$���t�sl���1[]70��3�n�����);�ə�lLaڻ�k{A���I�]�l 2�7�����w��^��^��JG�)�ck��t��rO\�r�Z�g�U6E\�a�\f^��|��ħ׉��v
</������ӗ���<���Sʠ�VE�#�6g�5�����b\0fT�mμ�g��\}��Ir�q�$p���2��\���y[�z�p�n��i���_�Mn��S��G{Y�YfrKY[����8�o���l�$�8C礞��6n{�	D��_)N#��a�� �E-�9��{�kE��żz�L�L���ͱA���i��D������J3R�9���a�;�ܒ.�A�'�~A��j4���H�H�j�$�ZZ��~KYp�*���eB��~��	������Jw�\H�Y�藹Ꚓ�7���ܟ���k=�!�c�z�.nRqa��/�}���wH���٥A��'U��r2�=?zܵ�^H���$lv>X�E��𠝇jU=�nFA�SfQ�����P��݂P��F��i�iQ7�$��G-�Ф��eK=l����!x�=W;v��犡\*���0C���$���Y���m}�/$L�K:��}���)�zGY�R]Lh�M^���|�IC�VO�Tk�@�].ڟ�lmD��995�DX_�����q�`�	���7;�إFd��r54prM(���4=����ُ+�:�:NI���1�M�Qm&�����tZvR���p�^X�?�+F�:��M��tW�l'-WMAӛO^��$�8�j)S9`���T�ow���ç��]�A`���&,p=�E__�y��kD3��̗��7Vw����
�:ސ�'|�B+��Ȋ�Y�<�f[��HeP�.�>��cS���^|^���0bR�����'�8cx	5��]WD����U�mE���)O,Q���]��S�3�nw`o�-���0SLB��;�L��`�֔��~���+,�k��묱5C�Zǚ��w��]�$�ZƑ�Ik��ǊRJw@��'��.�y�$/���-�'V��;�DL^�5���E/�z��G��]��蛥y����jbTJ6��9ꏶT�u8q|E{�#�u�E1bH�����0�w+�H4��+�w�����Sm���g���X=�T�<����{�ҫ�e�
\��M;�����ua��+�D8��1=�HT�$�SR�����u��O0�0T�mai�z3�nF�!@��gs"��dE'~���O��˴�g�]��!<^��U�Gg1�ϾG9�1���=(t�u��E�{�VU��̊"��>H�[����^hQ� ^�R^~�mo����iC�~��l!f1����'i�(�O�u]��F���U*�Bխ$s*W�JF�Cd�/��+�Ryam�����P@��)[�W"��3�5��V,��W�a��,����Ðm'��Uq���f]#�t>��lZ��8�,�r�I�����t�oO S�������[�<_�TtӚA#:Ό̗ݽ�{G]��mK7��� 6�'^Z6}y���y�c[b8�[��w���G��׃b��2u��__.�PF�O��Z�(b{�{>�`4�}��<�����ﶘ=���<�o��Ї�*(܅g}-8�C���� ���)1$��K%F*�rH���~��M5�7��U�G.��9w(:��x��6�O�)!�:��������>Mv0o,���3k����=�@�|=������åf�,u�*��xp����bnEd6%�e�:2q�����U�r']0���Y��lg� ��P|l{��Ҝ_w�b�3� �~d\���8�����\09��`���� x94���wl����b^"��7,:���w*����*Fn\NW�R?���&���}'����[�Οv�6���fkܘ2�E �wY����}ؓ
ZWz���,� �= Hβj��	v��qӊ����5�W)�����Bρ]�
2[R_7��2��/2���֟\^Ϥ�/	��ʙG!aba{B��(	�\�G��G�QH��t�K!�~_>��Y��!]<�Ξ�4y�k.��Gc%�g��y���c\�@��Cb{�%�;����	�`��j܋R)��#mZ�+z5���L��G:N������������C;��m���3���񡎇�� �?q2��ӃJ#����y�w���3�Y�(��ݼ���CH��h_�ӵ+-��ÖQ� ����EM����U{m��$j򚑠~S��{?�Ɗ"vv�ĩe%� /E�$gĆ I�4<^S柝��p��K����܈ټ�5h���=���泚+/��H��HP�9"�/q�!����y�g��s�R�a+�y
܋1<���q�DZob�;��s�=���gϐ)0�U�\z��aѾ��Q����=Y������a^��Z'P��W�/l��D@��C_)�}��<���{�lr�N�C�}J94�3Ox�F���s2W�"a�zKL?���YzT.sm���O	���2�穟����Vdjs����0����,Ϫt��q۬ǳ2>x6z7�/���G������9�f�-������_z�47�3ohv5�$�ʚRV{��l/�4!�ȆK���|�&l��X�	P��z��q��ú���d�8��cA��r���	� ��B�i�ӹ��G����ZP�P,O��xy5O����i8����>��aq�W���2v	\�"�+�	4��Rۇ4�^�U+BJ?`�Vt�8�{Ӕ����sWF5T"��<A��n��4�Ĵ�z:�w�᫪
��\�q�Յq%ro2>0�}���C��oC^a�Tae�t�\'�@0Iq�-�˕|��Ⴘ/���^D�t5Yp�T*�R��l�t)����I�梃~��N�V��j@o%�C�Lu'٥���v)4k> q�%`�UQٯ����r4~���GLY�O;��$�F���K���?٣������]]}��(x��Ĥ��>y4��h
ܮ���>��;rv�S��߾�7S�K n;�A!� �(����Ԫr�B%��̋�=�Yuh$�	npC��ݞ�$�9+`�Cf&�T<�+qTM�X�0 � ��3�y{ml\�R)�	�fķ��rI7΅���@��ڧ���x��q�W��%EG�T�}&�򦣾v�S�qZ�@��o+�f���<��KMg����/�L�Q*�~�����s�1b�����S�o'U"}q�ߡ�d����� ~���5�ĵ�䵃����YhJԳ�1:	+�h�ۙ2T�Ҳq��q��
��:���
�/�3n������Ѡ$�2��s�iW�y��GqB��i�����?����K�T�����,��
�鷦3��R��r"�d#��g5#d�Tz�m�ױQomZ���k��k|�����/�$)�Y���7i��Z����I˺H֮+���Q |�}d3�p?��4CL�V�[�>�r'�L8W��Y�g�b'��F����$�$�&��3�ҎM ԡ�Ƴ���ש�N��lI+i��������(��vi]�纙'�	d���)���\ ��zg����lg�s"��D�Z���N��o��˞+�ĺ
���$�t�O��~��*���_�b���O�_�hq���t��1���`��Z0	 ~8-(��9��-�	P~�'[��U�����h� �w�ł�3Ȗѭ8��0lf��̍���W�Q�	--k]9�����d���򱧽/�8!���G�$�[�	�&�m�]j���P�=���*sE�_mv��P�0�/�lT�����8���qm5��m~�ꕣ7�o����w9�Z��,"0n��_ ��HT4,�©����:�M�v�Hb6;�0���im[�� [O��X�cF�T!Y��y�(3����Y�	���U�@��K��}�>8N���1[S���oȪ�%/4H���h��9}�u]CķE�A+Z,w�< ��5ټh��Tg��fA����z�M�b-��u����|)�
�q�Okq���65�@K|$���i���i�F�O����|��O�U5��
�������Ј����F��9"]��VH�2>�h�d`��"j  ��˳Bb�*&���j/�m,��k����ĵ/3 ?{q��G��3&b��@������#��T@�\�*���4��Λ�\����xd_5��ب��p���[�R0ޤ��Qf�}�ps��T[>v#�@��>XyB��N������[�ǟ�NO�/y%1�,r7|o9KƱb��o֕�[!��C����Iu֙�Yx�~`G�=�\�!0kg;f6�#|���>�`�)�Z���`> j,,;fK�'� =TMF�4��_9m/�.M�%e,Xjm8��Dđ;�2���;)?%�!3�e�=_�w�
�1��J3,¼� �!���ѪXuA��~���)�v�!��Z��̏(d���*�xPGvF�Ʉʳ�`�pe��m;���w�6�C�O��6�����Ϻ!�Py��⾙ ��yA4G�c�2ׁ��HSG��ǲ��ٯ�C���<?5ġ�.�pw�����)�W���c�Ba�ڡ�}-i7\�U¨�u{�^�������#-�V4W�0����d8X�BeU���ǘ��{�T��ј |��";1Si���<n(���|=kJ��YnbI���XM2��J3n�d�C9�F�Z�P7��T֚��mZ}pJ	��h[��yA�� ��C	AxF�K����"]
��-\�4Mwe�)�5ǈ���p���6^������H�B�C�O����C��a�-�WheK�8W92�&T�mAtB�R���c��:�Fǜ�5p뇗G�=�q��W|i�'��@�Ӯ��"�9s58U(Id��S�����+��a�3�bl3�vS�X����09�-���6{�����PvK-A ���Ɨ��ǹs�a�j��q,����>́ ����u�X�����+����~���g$��y����s w#�����-����l�u���-ʇ�>���Ӻ���u���o{��� -a"����j�3"y�h���CI8p%Aw���˿L���?6a���mV��؝=�o<�)�7�� 2q����e:/n^�L��l�_�!��6���ڬ+��t��(m�,O��acB̀;�� �_��ԝ��X  ,[����A�YY�d%�rCdY��]M.0��b��R�������H�M!~��.a:�mTak����t3H�r�`�s�3�l�".Y�
{����h
�FiE��B���x�IH�2@���J4Z�&; �s��d�Jv�u�W�L��2�r���,Q[��c����(/�=>�m�����& �4Z�:�Lo�S�wf֫�)}?���������|�[0k�1]��jC@�o�ZU�&��O�~ۧ��NhF�~�p��u@����l4i���~^���2�V������HGZ=6
��Z�H��X��z���� W�OYE�ϛ�O�H��腡�=�"�S#��[�B*���n�79����1e��Rm3w+ �&��t���;hZ�(!��M[�[R�1j�\ �Ⱥj?�A���`v�n{�m�8��Ѝ<��V~|�~�j�t�Oj�O��}\�����Q���/�$�c��*?[�`yMg>;ёr��' �h��MW]ki)�¨�{7��s�]\�1�����P4����u	!��8{��5 v�-�Jm���li��Ȕ~��o�0D����G��������6��G?Om*�m�لu�c��Tڹ��n�\�M`kUY*ⷀ�;�`�<L��@�s��m@8m�v.��ǭ#�l�M����C<|���fbN��>t�yz<�S*{m�-9�N����0��jk�$���X9��J��q�?�C����tW��%h���w�
.�x�p�:���"d�f�^|���SA���ۨ�c�+�#��M�qJLS9bx�cǰ�]����3>��_6�!x��͓
nY!	�QO�:㷁���5�a�,�A�(%�_ZE�5�`/��r&wx0�@�P/��,z��Fo��-�d���^
p��rX���Qߐ2�v��xě8V�f�zz4�D��	Y��F0��4y�$֥!p�$6�>�?�F��	����G���\0��s�&���Q��^��L?V�V�h�Q�r8)�掽C��K�a��W�辽~z��6L��TJ)�ܬ���h�	�c��Zvh%�������>�*�١v9o_M""��:uOj\A6\��;5-�����ĂvkV
��N�uZ�\� �{7���� (VV��)��["������ya���u�g�q��V2;/���Ⱦ���)�Ȥ�y΄b}n6I�����)x��Λ>�~ㄧ�.���E�/N���L�?�"�ċm��[^fv�ٟ3�U�\tsNIE��	�ev�l;1H�S6��1���.C,���v���V}���D�	$z9P�ia��{Qz8�(Qߓ<c����1�qK>�R}�U.��#��&�'4� _/4��;q�𢒦�»�0�l&� �5��[�,W�Ǽ/ɐ��
�w	nK�__�eD�
 ��%߼̋[HGW'{�O��ힳ��?_������?;�f�|V�qz;�n� <Y�+��j����a;�R�U�ך~I�
�����́8�cb�%[��0�������C�c+
Mdf�����0+�q���ًk�������=�	!Ow9�L���r�	&c�L�xN�؟��|W��}��nFIi��˛;Q�L�XJy����I<e7Č8��w��>�n�b���i�	���Z���yE���xK�T�P��}�|)xgJi�유�w`��ԣ�@��egz�)������è���j��(}1��������Ex�j!5�#���V�U�e�t$7+���Ugm�c�I��x��U�RxL0�j�W6׍�'�z|qA=��!9�5gV���72#�Tc��Z��b��~��#!&JUO�kEe�36�:�1��M��'cְ2oqd��QX �O¨cV���z\�N���b_Լk�T�?�j�r�<�6�ө?��Ouf����=� ���m�Q$���b#�������1�2%���V䰩��u�i�-*�p����U�O��F#��%�6�^������C%h���,�g5θ���C���5�+�qd�q1�hHɂ��
*Hr�C������F8��<�9WG��y���*N�)ťszh�ͳc��c���ގ�h�
;�J��uc��az�<���	R�i:����Ϋ��}�7�ܫ�*ɪQ���|��p9��B<"8L}T,
�9�מ����/���=����L%��S+�j�RM��F~�%R}p�&%�j�����_�}��Ɉ��*��jAe�hwJ��¦l&�c���e��<�����?!fN��Әꖽ��1�:�= X��Ȯ��R�Sfl�6f�jh���c3-��͌&�����aF7��0k`4:�gY�9�P��"��.�7��N��>sd,����m���)�z���-p�bCbV�1*sd"�Q^�x�04�~vw��U��ެ+L�6����e/�� v3��J�O�� �w�d��Q�%��[䘰�#����X<��dL'�8n��0��s�ۘ��}�S��W���u��_e�ʛS!2�o��dt��MwT�q��v{?�����;$�!	ZWt�����~�!��8|�I�M���<r�\a�#��&�����S+ӓ{�q�^>_���e�Z��kiu��Y ��Aa�VRg>�b�#&���p����j,)�b��y��4�EPS��v&�C�ڱt!��G�鏑�tO���Ɂ�ʐR�L1յ�+D?[�͓��b���i�Y*4Wf2���6qۻ���c�""�B��
^B��n	hZv��ɵ�H[�%��Lʇ�R�B7����k�8�R��DL8Sq�8�����wkm�[�y���/����ͷm1e�
�)�8��9?�<Mq]W�5[==Ȣ�1���K&�$4@�dm�{�;`_�%�%Чh��x�>I��o��ްX 6�Pr���y��������5Ѷ�]�U�A*V�hc\��:έ3���o�e�)n=Z����3��()����2ObT��sB�l6
ب���˟�K��3O0��kä�4B"�*eY/L�}�{��X�<��G��v5Mt���;��������׉��̡d�<�\�<왽89Z��^g~ҩ�7����@�ׁT�f� �.�5`9�VbW[X;ssz�ei-�<�V�uaXb��?�s3U�NVk:ح�\A�汧r���� B��-@�-3��0Z'>	BM
v5�q�_c�7.(W�{*�}+H�
�Q�ʈ�v��Z���FܤvR�#�_�L�aB��%�+y��V����R�A���0n�`���Ot���;�B�{�hv�NU�d���|��$P���ʤ>�Q�&����?�[|F�'e��Nb�żi>|ߘ��"A>c����^!��&^�H��4��ľ<z�y>HS�)�z�s#Ő�Xx���hkm^����+u҆����%a�r�I��F$ҭ�x�`�Lk���\6�u��6hm��^*rʱ���Fc��|��;9vn�# ���R�):R�i�fJ�kr;��&�8d3�5$���F�|���p�!+j�L���\� ��t����1>RI�3�1���	�LA;F�4����i�J�?�5���<5�d�
������?��C��4�
�Dr�L~�9H���R P���h���_K��g�'����J\�*q�� ����"Ԁ쾢wzUyˮ�?kmW���F��%�:MU�l�ĥ�����`z��	��P����8�1��j�;Cʿ��XR[��6�؄�Z�hw�X+�|Ğm?��҇�n wI��*{�d��2C�Qy�	,h>q0�gi��� �7��/�u��i���w�-3)B��L���6�N�U�uCR*�15��sO�3A�';�G�~���&J)��D#�ɋ��4vE�Ͷ8d �-i���Xr�т 6>�o�uv�-�716}���dw�@8Gk狍z�_�l�,��W)w��!%XM���QLl��k��)��L=L�Ƥ�5,��A�4��K٠4v1v�6n��B��m;G��K�r�dFH���>"��F gfM��~ϢQ��w69���\T���&�}��z��9 ���K��C��>�G�r�s�`(m��l���hW6"���/�t\�.H�*gk��	pqx����������0X���w��:�]ŪL���� ��#yiM��Z�6� R_{��FW���N��*>�xIF�}A��Ӥ���N}3W^��)�:ڳߝ���MD%����r}�!�Jv��#�7%����2!l��>.�t��� �/������	@��_��M�y h��@�c��	���� ��R�~kÄ�2���ZK{-�W�O�Hn�*�c�ӾM����<;��*��2H�0 si_��RH�����7V���;�oʕߚ�I㑙{�m�i�<������<�=���
(^�\Û��vp���!�����a߀��5er���u� ܡ`��������k���Һ#H'�5����A�@d�������2:~"%�:0�@���t�>���\ڞ�%�ǹ���|
�3��3�Ş��mڄ�!)Q�x�ʏk����G� ���I��L����m�؞�����mk������O����/~�"�n�$c5�
ȃP8��1���0-��.��Ϝ�"'��|�X�]U��Yg�'�,� {;)T�$��bk2��QW�w�rN�EZ/�����c�S�r4�LM���%�>�ԲVm�^2sNďt��e�_r���лE�;�UR�&P��6P�qR�e�N��ma�5Z��%X�D�� )����k[ W�b�e�����$����:Ĩژ�X6��`���C�#h�pp����ec�?�� ���%�?��?���s���fƐU�\=�4QQp~'������"u�yG��iy����&U�s8�x�Ј�._�� [��x�e��<�z����1<�l�Y�6d%���$C����f�o�	������/��E�Fv�L�#N�����$k<�d4@^�z ��AJ�8J'[!냶��0t~U�Fs��$ݪ~�������:h�ؽ�K���[-����č*a�DE��P�ˆ��5��+��[���\j�::����AH���RP�.ǐﲄꗅB#uy
���#L�����>���0�
�̤i>Feqr���$��[L��R���������B�gs��K:ot���~>Ӑ�װK�CGY��`�dr)��D�B�Q_3qh&±[��6NE,G�j�"5�B�ڒ��.D�Y�+<�vOoEN:8�@A�	$q�P�pUu�U�>��vP@AKD���\bx���C��g�jnT�w���u�,�$:S\���m��G���1���/7�L?�D���_�)���W��6�f�㇕a���n2�m��2ғ��F:۩ɯ�`@��L�090�F�/��|�8�^j8GF!�����N����ʝ:�X�~j��h�9��Y��ujr�uH^C���o�Ţ�J�e��VA%��ڔ`�g�#F��TT�����!��pH�4�h�M8����M�B�{�����"�̯��2�]d��H,{kV�X���V@�����N�:���O�X7�x. ��e&��<QN�
�\K��1�������EG���M�mV�ĭdz�� ҌAcb�0��P?nJj��K����}�H�8X���7Nv-��kC}biU���Z�k��)��x{��=�T6�V
����q�gq�+ĕ�i����u�����#��g{�Ր�$R�!�gDe��E��\�.�� ��T���׿�s��/���<|w �z K��ղ��3��^V�&˓�D��ud���8ZP�&���	��_s�:��^�1�6�4�h�b/Mr�����)9�T3����P�X�F�}���&J�ee�2��D͹��/oV���j�K�����F�]UsFkJRGX��e>1���-�L:�ī~gx�	U<�HB�6�&����������������3�c?��7e���b����g��C�I]��嬪΢�%߀D���J��f\��Za�b'�5�8Ǽ��KҊ�Ҽk	�N �'.-��!N��_����h�U�k�vD����[�A�yG�؂Z����q� ����ע:�ZP�#K��v����ܱQb�O���l���Qyp\Z玵Z�l��7��Y��� �0������䲐mZ�n����͢���J>Fq�	��˸�# w�����M�ў��⿙�6��UO�F"k�y>h���~�7'`K�	�:_�;*12[�*�J�wYRt��\�|xLFl쿋`c���4X "�}�����îO�ѵ�0�k�ubQ�z��?
�.�F"��M�T4&!�N�;Yz���mi!A|/����N�]�qx�����x=$��*��� B����<� �8g���΋d�	�_����,�c薴��n�-꺌�"����-	=�p8Q��A����s����u�Y���I!T@�5�l+@(���z2l0B���Z5^<'$��I�lh�?�=�b�J�<�^.]9zW-����h����	�4b_ ���P�ǚn�}j�e�du�(�J���Z��������_I���L�/O?tg�(n��N��D5�z閘:	"b�%s�ڒ�����Pr�����3|uG'�����Y�Dy�
-ٶ��0s�!m�)*轄=8�F�2g��}��W��vFQ� =��{�p���$����;œ��O��b��x�D�M���[��Bg|Ԡ��r}�S��#ee��OĮ��6!�^�;�cJהy]H���=R���b�q� L��?v~�EI$���Ǩ���-V���@w2\�mM��=�C�Y�r�?Gk;�� @n�H	����	��ǴqKӌ���~����w}��,�]�h����%s4�!��|/�~��n�#mk�'�r�-}�O�W%��՞��v�Vd��l��/���"oP�5�i��u�BP�/��'}��Z0�8���`;iz�N���������<x�H̗z�ǧS�P���t͇����@'�|��A�l���RX����Φ��Lv�v)�lZ��Sa"���e�6~Î�[��g�Z>����A��#���Wu���L�RE��	ó���t@�Y9���7��rDps��C:0����]�\�J=ٿ����_��x�A C՛�_]`f�(_��1��7��w�GkI��㤼��^�v~���7}�ܢc�fIͻ(�h�űU��Wz�i)��R$��i������V�:`^�Аp��~�uS��Un�BJLe�]Y G�&��p4�������6���q��5q-=��u=��!ԨҞwU΢��� J�m5��+��ZpG�PkЀH�F�ffn�n;�ׄH�tk�����q8���f��)���)�;>Hp��{À �u6z�K�xY�u}�z�*R�~;�6������>y8���1O�ev���*��?�2�e]\��K
�x��`�Q	-��<$��ݰ���b�h�=wx���쬇��0т摊&��/Adb4�<���+���T,C[���~����Nz
�L4@��ɣ'�~������ʖMLD�d�|Cf�S��Y���N�v�O�N�QL\��9�{����Zd��[V�'h����.L.=�o
��֏���B�X��i/��T���h�@[�����T�Z]��R���Z�2��}�p�Z/254�0����4��h��;�έ�V�;%)7��ř��ܜ���Ok!i�a
�&�͝)�;��4����a4��@���\h�����eo쥦��~�,.��<�,0g/ρ��(��[����.�2��P2K���*��u���{ �M��v���'��.22�Z�"��(�s�{o�-�L��r�X�bt�v8f��TFPM�~G�ײ�}��өN�����h�`|��㣀K�~��'oͼ����I��`:bnZv���5u�x�[�.f�_㯺+/�쀅��������`Z�/��{���];,*,�?��G�Q�Zʟ|0	�9Զ�N �6z�8>IH�jD�:FF���U��ࠦ�H;���������^�ir�{�9@$:��-t�O}������B�kk���Ć3��Y�j�L`�#-q����UU5�"c�ޫ4�)�\�9@���%8�/3�����7g�o<�^~u���f��
2������|[f��2d�~�ʶ�[����p�0{9��{Vw�?` �3Zh�t�^|xy�|n��AOy5U�����٘�ٹ&f��dc��~���s��I��8��R�����3��hG�F�8FI�V���J�� �8D�NX�6.� u�p����0��ݒZ���m�џ���)����i�⹪�w�q�at/i�D��j^-w,F��By\�".W��t$H��-��EK$u���0 "2����3=���\{�ʊ����V5g
��==Z��;$�VO�p�D�NǶd:
/q�Kѿ��*��{�@͵`%�@��� 3m�\�$)
��#�[���]di�S
��!*U	��ӹU�W^c���=N/���)����>(9-Bv{E6c��k�f��r9�7��sR%6B���x1��8m(�/E��fe{��HùQ�٠s��81P!Oω�v2�|�,U��UѨ�e_�P�s�(�#'$����#�(��2o��7�6�b's�9��m�`Q�`+'��R�r=z���*���f!TNٓ $+�!Ҭ��1��K��%��,�9�cE���ŕ����T[�t�=f�P���E���q��p�W�Q��۞�=~s^D� [VP� �V����B�©�`� }��M�2�Ȝb��%��vu6�m��p����k�-��Rh\q�.�|��)��P���5Ӓ�"_(*:o�UI�����T��v��P>m��~z��*��VV\�����]�⏂:�� �:��e�hbΧȣ��t�=���u�����UW��My�K��הt�sj�����FL�寷���R�c��i��H*�(,z��e�nAz�^�b��1'M�Z�0��EY1Ƈ4)/�n���/�Q�6��W�����ɯ� -���B̵^p#�h��H�"�-��-#��9�mrC�zP�aA�/��<�ϽTZ�k�	�����
Ѽ�X_�q���IT$/+ȁ'�?6@\��P��e�s���w�u(���ME39�Fd4d���%�"-U����J ל� pAJ������d�+�[�xe�e�`|f���xn���
���'=s&T`�P���-�ӻ���]�3*�i��I�#:sET�����[��n�K-��7"�����e��`G�� aN�Ǝo�D�6�|H��s�W�˷� �O�Y� ��`�
IёD���E0��R�6#M(�"�a5J�R��OM9��MX�=3�<���{+Y�ٳ�>� ��;�8ቝ�:�a�Y\Q�+�����"�x��G��	un�'�%Q,���X)e7r��⮆$�:��J�M����8c��7HCLjb�!YOMX���|�$��<���$VqQ�K��}��	�ފ�7�����ϴ��P�P��$�fe�ƺ��#�ٱv �N�8�[&B3^�f�@��b�H ���F��vͰ��ߪR��]DHm�~w7��RA(�y��1� �ƚ�@�X3K�Ѫ4�Oԣ�Z�|"��ۉ��_0e�П���ޥ��wq�9$I��CtN�l��0t`��⤓�Y��������`�N�
8wH�c�2�����m��;��d^[d碫$�N���5��W;�&:k�����՚���� ��R�4�7V����>R46� GX��b [s�*�>&�F�3�X��O�#���}D7�����v��Tw~���[�u���~�C�+����!	4�%Ű���:��blݎȁ)=�
�E���{ 2fGxY�5�}�0������V��3�@��&�_m���y��j�=�΂���x�����;�D�ْ+7�;��U��/�r�܁q*�������C���m�e'l�¬�
P��xV,+9ZR�:_�/ep��lו�'N�c�%Z?�O���,p��#;�H]3��i��#�N`p�D��P�Ah4^S[�d�����z6M�o��s^m�X�Ľ!9����2�|�V9�i�:)��ea��7�L�U�My+�h����:ɩ�����-�	�ui0I���2�p�AS_`��`�p���=&��=L>H�xs�[�!��)ꡱ2}���8�� �D��ǐT	���z>6���}$O�؄��k��y��ˮ@�[�Qf�H\\��|2��S)ۮ
�a.�������]����j*�n�Goz�� X���V&�l�_U~9������Q���
�I^*d�g�̂��G�tR����w7#�wE=�x�Z���F��bI����{o%Hz����m���Y��I� �^����� � �گ�.�smo4���P���氣�������U��@;��,OA� ��Yr/K�J�yJH>[�����l�*���^�/�%^�Ù�$Àm��y:����m(D��N+Z:���Ɗ>+���#���N@m���V�X��9��Y)�C,�y��߱  |5n(9�Z`��J��A��&��bo��d@<�4:�Pi�"1�C|�+b�����|�1e�E�B�����d����:p���%�Ï�Lf3<d>�V�ܯ���Db�pQ�:%B*t|�҅����9�V�7�wT�NI����[�\�����R�o�n��5yk�b�T�l�9�R#���a�`!Y������Q�{}fS����適��|�7]�%��1����a��7�������<���N�V��Z�l ��*bS�"\MJ�ٌmA�d�\F�؜�@:�B"��PSyjuo�	y�����OY�'<QF�ɂ,��f�������G~aA�@��?�z���?鋔m�b^��#��cc��}:���,�h�N�ow��^��g7�� ~x˛��wJ7��eh{�:[���DR�&�\���fP��:�1�S�I�6��v��š����C
s �1#x�JYn`�%���guc�g`5���[�썑�v�1���4����[�
nW��( ׯ�XD�'��ߚ�.���m�4�;�����C��6X�H�J+�i_&���@�%i�������!��� á���I���[�nQnw��ƆMS��p��7��dڎʹ�C�����sj��<u��263��g �\�
�)^�v_x8P���"�ף.�K<,�zT۲l{\�����ͧ�h����Ip��qï�8�SF<� i��k�m��n)wn��i�~�ӈ5ZYki�P����MR	<gM�n)&�'�v~X��׻ ���-��fU�3�{F�b��Ƞ��R�i��3s�L�g��n������|~
�Jp0�[�}�S�;����"A�]>th�yX����U=02b'JN§;��y,S��7̇������>�?)k�M��G�2so�0,���]�&Tx�(S��I�h�m�������@��{=5�p�M�V��e{�S1��+> &�z��6X.�����+���a�%6�I`�e��Г%N��s}���ơ�k.f�@�hE�ڌ�s5�?0�]��'��@ͯ�?F_Q]9�>���{!o}Vɦˉ�P26�"��g0Z "_������w�>�f���sF�~^�^{V�烸%��{^�(���x_�����Iu��ww��IȱzL!������N�sP^F�*�t� �/� C8a �c������~��q;��� ]��Z�-EqF�ˍ*-әP%,嶥�0�Y�3_m'��&?"���N(X&0��?̓W)���ק��T�@~�P=���1��"�Ɔ�i�-h	��%c�=�Ƭ�Y��4�?����@���=���� b
�G�u�����m���a�	��0�ia�E7�������ml׊D9�m*�,'����5� ����y�}�z��ǁ�������u9�,h�8B<�����Eo�3(%Ơ����Q�f����pB���}��e p�٭*+��
#5�r\�jn�U�`@�	3UN.�̜d�GMlTK��a��r�o�2�_�>x��o>9b[�N-�`0�Đg!�}.��� "t�e?ߙ�͛��B�uG�1����'*ҥ�i��\晴 y�>S?U���h�@�Ξ)L��b|�*��g�Z��%N��E��P��g�kY.r���������D�s����Ob����̲E�j�^�7��>j���V����'�?�)ђ���@��M���z�Gs�'i����'<|Q�d�t�&�{� ��0�Y�q��>"�?$�6\d����8஼f:����oĪ������_��ڻ��]�	h�U�H���E�$�H,e�����VH��
�x���%]���<1~Ikh��-�S�_7�Hk���ITS�6���&%�2!����C��b�	����w��7�&܎�xr��O	����סL�����v�K�"�g{q���3�����L KI�]z&E~�S��+�E�߬��h�3v�V���jڸ�X�6����o��s� ��Y=M���;Qd2-��CT���Z�8�:�FAWd�&��{\�Hyo\��\?�:�W�:�6jQ��j��	�D{rH+_�+⴦�E���ꝹD�m��t�a�%e����� 護5���N=�I:�#�J�#FZ&2��CRW� �K&(�G8»gn��7���Ʃ�7|���OX�i�g���4��!	f�O���BĹDX|�ׇ�:zǘ~2��M��H�>qU.��n�(����-�li�����b2�����N��dG(���E�n��r��_]E3Ev�����<�O���u�"L�
�:Cf���A�r���!��#�p%���Y�4���Qr�F6�S�q�w�U�Wq
�/����lX��P��$k��7�B*�m�3�exh	�m�X��m\����,ы`t2���ɰ3�]�s��Z��.\��+@�z��Ϲ�Ș��*�0ȭ�Iؽ>�Gɮ��H�x�v�Jl�F�0�s�"�� ��\�u�C�!i��R�+�^�p������ΣX 4�T(���\�x����G�E.:~	�������vKן��~��i.�ʏ!��(�1������`����@�hj�{6Jt+rѩ� Dy7�.�[�@W
U'I�D�lHDҟQ?�l�0��y|F(����@����|�L��uj@�G����3"c��1�/���-��|�|���&��Jd�\��1����m���G��ڠK�>�7��=�v��y��'F@������U�g��h��.�B`�%!����m�BUW+A^���$�fa$O�E�)�[8N�R%ࠬ�,֩��PN�v�;���c=<@�w���p8Z� �0>Q��du���gI�(��~�p��e4� �?�`�}~Ǝ�SVqf��5b�:l.%ю�'ˮrЭ�>>�yC���{��ν�4�"�sX��i�M��kp ��IĖ��c&�$��=�X������_Q~N�u τG_�$L��$�2�4(�9�2���(�s��(�T��l͊�+����mL�u)T,�H���e��jGTN�q�l���#�G� ����$�X��w�G� ��.#F|��~��>��+�3 ea+ƃ�.�nP���˶�)#@yyo]��_�K$�jW�s�'���1�U���> �0���r�S���2�*���#S��Re��1�� �����:���|��`��p�UQzQ05�~��0`C Ӗ�W�o�#%J �n�w�be{���!%����/����1D:f���u��(x�?�: 2�r�]�-W���a�ye�3ksE���N\
��@/�ɸI���3�!Ź˿y�b��	�;�^B���f��X��|38
-���s�M�"TrJ��o����S�ׅ'����O��鋘���>q#ҁ�ؐ���-�t�gPu�^Nf�	pO��k� �����ʍ�´A�ѥ$�)��HQ��ǘC\����ڊ��18y��@�Ienވ%'?���A׿m��d��37�OA�VD��=���������(�)^�2*.4lY-ճ�L��� Y�y��^��7����g��tT�x7
N�/i��7��2�t��_f��c�"�������:�4����j��z�|r��=��@)�S��fz2H�UZ+ںp<��;aN"��̩+��ܗ�"q�Xm~Ó��!A���q{ h%v�Z+�߄��7�69�`�|��HY�#�U����{Lgˀ(}���om[�B��
�W��C�мv\-`�(e͛7��&zx��G���g��|�'Qq�L(������]�	�����5�����E�[lW��6X%�A���/�h:�_���B�-�G���t���G�W�}n�x�ؓ����������iK����wv�M���?�ss��L�v�˺�9盡��
��&���{��8�<�����]��(͕�e]p���4\�M�:XA}�k1�/�5�~�Az��f�tig��H��,g�c0}��t#�������$SȻ�P7E&��[��VY�
��վ
�݀z���i)�1��j� ψ?���d
�R�1�\Z�����P�Y��~\�LjR�q�ni�+���#���F*tJW��y���T�L`��?f6��) ��Y��J�y�~��#B��ÕT�$ts�Q��������l�Z$��7�s[�&-�$���V�B�c/!,EQ ��a�����=��=(�ݗ^S(��({�0��-�"�U�����_e�^�Z�d��������,��5seH_�'�(Gb-{�E����%���mpAh'��V��?1�V�5��Q��%01��y��xO��-��K �+��M��Z�+0���(��-���V+�������t�h�CM�,E�t�u�hXUx5�)��g�@mw[+|M��9���б�]s�B�l���>p�����R��uC��؜0�ri��M��c��H�vy�V�($�)e�:�{GSkN������S����B�[4l�ЦCv��_�u��������9����Q��Y�	���?u�|Ӊ%m5�N���aա�k^Ș��b��SmD���C��Z+�o�#M��R��Q��Ƅn��<��&�j��G� ���B#x��B�J�s��)�@�{���Qk�T�ǳ.���C���?�!�D1���0� ���aHn��E��,�i��I� ����oag�T���6���;�x��a�MI:�zZ6�(	����i���#�ŉ������߸"ɜ��}�U4Ԁ�$֊��n4��I�����Y.����=��O]�R�#!�ڦ�0Q(*�;չGw�S%��P��>�{�@z�Y��Q�$XpD@
�ao�ctBV����U�s�ƨw���HMJ��>'������P��ni��VV�t�O�c�~*> �1Lh׭��F%`�Z�� C�)ɒo:�5��Ȅ�!*�e��d����뾩��f?��D2�����	�T���@o��n�g�+��6���?W�8��9��'KG���
:���ܥ�x��F�1	LF�Y�4j�6U�*wƐ`��i^�)'���5ŗ$YUDk��Fu*�;�%-~O�R��jji��{K{���`�%�$"� .�]ncvy`WZh���m����z���2������R��n4�B<���Ŏ��cN�$�4��H����q8�ز�/@��?���B�YƠGB
8U>w�(����A���me|)d��
�:q��g�J�M�򺛭&��l�F��Ҷ��:�vξI�.mh&���l�����-vO���L<�A;`�)�l���
x���I����&`��MΌf^\�O�F^�F�6p���iv�q)Nܚ��2[��L8y�������>G��Z3��ϳ�S�DAl@%����)g3Bs7׏f��m�#u���`[�ΪCn��~�����rVU����ĺ$�h�����Wh�ϦZ�L�S��W w���`:��p�`移��ݒ�b�����CV�Ta'+8 ,J��5�Ge��B���:^1����*z{;�~��q���O�F���sj[Y��}0Cw>��\/�P����]��aT�]T��kFnw�<���3�Y+bu	�����&R�|
�@��C�ŏ��hIGt�_{x��M�U����=l?i@�X�b�H���?2_^�/�:&����=S��'�'tCWH��Ci��^���<�X� <����|�6(��Z��t�f��t�zЂ	xH�y?�#t�S��s(�op��CTQ$H��X�_�q ����'}����,<b|S�+��T��T����9�Ѐ���U�G��G�ՐW���Iij�ٲz�R��n,�P��\n�!�q^&�w1���B+o��Y�D.R���ٱ���v��a�k���W��
�I�u��!��Oq�����+���^T�	Y��� 9�9���C�p�KtTP4�Wס,�@,�����ث��sl�T�Pgs�+�5L��)&l�U~ᘌ�]�gB�(�%���?��?�6|@H�1<���rY��f���P����D����	$ǽ�69�QMS�dV��e��-��V�a%��BAL�#z����x���/9Ӓ�B71a��j}�|်����[r��3-�a��WQn�D�f#�t�{�� �ϡ���ç��u9Q�U�I�MR�a�{cy�Ύ��h�YQ���	*pփPw��K=�E�U�0����ߔ|$�=ᤪ����&�4�������L~���;�Q���ʸ�T�1���!D�y�>?w�Q�"G�u��5�*��]���	U��X��xZ:!�+'k��m/��}]CR�����1l��}���o,k<�j����9��r��\�\��JnIՉ��5}�>y.�y}����]ښ�!�4��kz%u:5�-�٢Ś�8W�	ޞ$�V.�N~Q��sۺ5=�q��Ҷlt�����L;�Pj�ߚ�4�����{��@9��	(qP�1:m�,R{t�W�=���K��	g)~g�Q�J�!������:�ڒC/�Y ÷�]�ӧx�S	�B���~�r����u����5�V��4]	Bz�6���;kaT8,bk@�@� q��59#;z���JVW8'I�P��yj�{H&�8!z���N����K1rz^0�˦��1��?���ͩD/�)%����Бt��Ja�j<��˷0����YaY�Ҧ���w/�[wj�����A���h�{BI�N��F���{�"wvY�³�>����
�x� F:l��O胜M�A�:�oJ� ��gd�������$��M�j=�f}3��u=t(;��g̔2�2���e`%��(&�:j5�
iWP�����aH<X��}�g�_~q��Z�<uۅ>/�2n+yP�Bt	��� �X���0s6�t���`�)�dY��*��e���X���j�!�1ްu��V�qA]�*&��;DM�1??�iwNG��U!GǺ9�A��ԗ���[���	B�CG�\�W�� �c�_�ԛRc�/��o�O21�@4#��1:HŶ�]��Rp�}��H�xR�Z�^��s���zg��2��K?��؜�@t��~hb��J�;������}b���8�0�P^�M�����gyQ]���<,�El�"w�]�W�3�#���E�LK.�������w�8B��"]���@"Q�h.�uz��XE=�ݾ���̍��7��͹W��*Q�OݠϺ%k�¡Zr\���F�����^"VB�N�G!�z�lZ���.dݜ�5 �Us��s0�u�b�~V��ą}�A�[LN=���u3�G�5G�J��8��*��>�k���Y�f���Qn�f�A�N�g �ȏ���X�(���tH7�� c�@�9��$��(�!#L�"�� �֦gs!D�f��RAh�&U�U8A\c�!��13�s�bKc�;��{ �XX�RufǭC�̀��n��(�F
A9r���#�� ނB�v#<Z+��R�˯�s��Nbn�YF�����9���=Cp�p'u�A��u^�{�[�uL=�$���9�2b��r�@��� �<caN����_-C��P���e�k�WfIב��aU�ܔ �tD�'�R��Z�����2��m�O�����l>�WI1���
��ۭ�T���3��'��U��)�AJ��D+,�(y7���ۭ$���[[�k��>�ts���3�K�~�У���(��phCq)�I�rbf�w<��b�`m��*�O��Y�b61(;��x�T��x�f��X{Y�L;��P��$�g_}$�rVI��R�����$_T �gv٨�v�^�iG	-�>cp�79�Z�ѩ�$�wz�*I��G�eN�Kf�a75'�=���H	G[���H4�)O2�,�b���N�?w���/֐�2r0h#�=���n�'�X6n-�X�~��C�_�sN�'��$&���j!���ُYͤ��T���1<Ղs־0v;S
3bB�N�5{���G�Rb�=D#��`cr"��m0Hh����Q��)}�Н��ߜ	t��������Q��6G�����h何�Ԟ@�mO����\�_��t[��u1���(`�e�̝�^�Z�k���# 0�q�h�����g�e�'��։٠��U��8�aJO�.&�@�j:ף*��&�T��Tu�2�$����^Л�D1��`Fie�N-��8?w��wF���I���"m�u��]�{NFl^�1������W�è���h�����^a0��)N����1��8-t_��7�)���'�0�k�Y߱�mSk Õ`1�uJT��%/Ds�l),�[�����\n���G_�r��e���͞������I�V\Zdy��d�4�1�\%�阮�3�lC�ew7�w�k.z��Y��H�Ģ|�1�S�}U�%��8*��6��a%���";�х;�3�7�)�۹����X��ق�*�F�Q�������p펶&��Z����>|1���OA�&�"U�b7���IH^�)�V�d�!�$Rc�K8k��c��D��Sֵ�ռ�W�����l%�6�sg=��5��X�@rr�9�A�#�B��A�n��JԵ�M-�$c'H�V��|��`f5��$�^'XBF�Jp�j�XN�����W�_�c�_fxn1�j���n�β�a��g9��*��K�U�E4l�(Ő�'.��;Zն��NѢ|�1��ۆ���玵��$~��oW[(�xk#*X���,����r���֣����9&�����n�O�%��>��\�UYI�B��l���VᲞ+�%H�_f�<	��7{�_M1�0��|Dt��W��;xdF����<�U
�O�}U����b�z�5G�F�W�{m�<�	r�k�X�o�H(�@�k�V����|�ݩ��c�G�ܻL >�%��6s���񼟮ך�(�rY�A�8`��	�E+Us�y�Ƀ���R+�5���h��}�Dl×���u �x�l��Jd\��{{�(���+�]`�7��y#S�v�jv�X�Ǫ��o�PqU���ٛ����Nn�D9)R��FE��#S�m�!b����� �,$�%�Z����L�y��s�����c0�>?��pMo����Eԛ������|%JQΰh���&؍��-Q����ki���N٩Π� �6g�A�EJB"�o+���-�žcK*��X�6=���/E�z�Im��\�6�]��j��A���Q�T{��r4��O.~	zo��n0�$��K�t<yynF�݌�!��
�X�������X���Ə�9G\���e��NXةѨ5Z(Eb^!�@�>d�=\p]g������*�O�4����E��4<lU/��T��m:2��
`����E��E��G�2�D�>G���5�A�t_�EN�q�)�[q�L���M
�o���!SrZ���ݺ4�`��yu�Q���3נ¥�[x+�-�k���P��+��I�,��a�f�W�=�#�)`bl����sA�y�|{r�'���/��Ѩ��f�s<���T�(\���KVD�3Wi�s�"Q[��3{��BLu�(�L�#[_�uƎ�N$��b��{3��Zye�dTz�W���t<���{���jQ7�f*K�o���[<��e��qA�T�s-.�Х���e'�w0p�֪'�}ظf,	]�.���ۊ<p���	�����~����n��6Z�Q��?j��#bSh�:O�Z �F~T���#�[�t��qX���	&�D�d�<�F-��ѬM_���R��z��AN�*����/VA���:+�w���M��|s�i���ҋ���ǻ�&qY]Ax1�i��o~"}������m���C).����Ҙ�Av�)aMY��9*N��x%7�����GT�� �
�#d�)��h��?��[�G�Г�ߩ+�,�a��n�E�w��z�w���(2Kt���*�)�`����a`��JY	���F��������Z��w�oP�L���������O��
����+��R>��g3�/,Duj2��YC�1����W��E�9��Ǌ����!ҤA��+����GT�	 �P闋p5�"�ͪ� �����l�z�Dd�.�dS �`aV�~xpp��BËLn�g���>��i�JNN��XL18f�odH@��=n5�%6�l;C��Sq�-J ȱ�U̘&�y���v��aP
;]�[��DP�w�.�%gNx��l5^���|ˡj��Y @��VJ�Z�&-Ę\��b,�/�S���p>	��0|�8�v�M���K�E�B.�Ʃ@n�)B^C�d)�������5�4s��?y0�`��kH�p�ј��ː��'��<�vg��}�ʀ0�<�ј���	�I@�q��3�N�Ӛ�
���.�=��F�_��=�u��T�b(Yx�8�Wz5U{�ϟtw+���>D�V��f5;{LQ�S85=n��؈k�󉟔�����4�9c&I���-HK�����d�sw ��2���+a���}��@hǫ��^0�q}��ׅVS*���4�%f���Ks��X���$�XB`��I8؉J��$OF�?�{��m1������&�a��tf}���I�j�q����+{֬�K���MU(��⺣�>��W|�[B~F�J���6Ee|G�9���-ѿ��İ���Ԃ��ޝ_���B	mA��B��M1w����C�0��r'ws��',\�,�F�'ȩ_���z�[�vٝp��~oBJCXS�RUI�$�Xg�]m3�Yv/L'������z��������}n�iJ��!�0�H
�K�u��7���֗����f��$lv��Ѡ;Z�(���Ưɡg!��]|���`Ğ�vL1zŝ� 3{��=�u������GHq�	��!� (�Z�����A��h�"���vr��_H�BAF,�>�ģV���c���#�>��V�}�hf���ŕ-}@<a\�7�H��A��� l�-6��5��Vm0�'hVF^0���4����Z�+ԞN� ����w�^>��j�y]'���mV?�4"I"K���?ڶ�����Ų!O�q�n�E�'�SN�n���K�
����T�I�w�z4Ê��P��]����i����<M�&�C!�vM���`0:LXi���~*W���j�ͧ����u�O���km4�a�-�o�r^Yg9�|��1�stp�L����@�ǄN������vT�V� ���@F�|��&�7>�S��	ha['5����r����RKE��ê�=��s �y����s�A�ˑ�p���|=h�(j����)}1x.�l�Kқ�9ڨ��11�ޒG��.B�+�8�nǮ����hr3�B�]��-M�v��(��S/�q�F��oS���L��Y#�d@�Q
�n /�Țq7������wnǗt銃��+��~,�ѵ���o���^PN3����\<t	U^PV��:#m>[�m5�C0������N�S��cس�a/Pr/�(��b
������������;��6.����-��q�GFn��'��j���Q���o7�io���Gب�������,��cD4�Fm*d�ǒ��$>(��Sh�{3 ��[���C5�b?�~����X���	���e���^S7�b�wϵӺ	��۽���:��>ZS�y�k�`��K��kb/��-�dY����B�������j�%g�m�����r��`F䚐�3�'�V~G|Y܄RI=��=�k�k�y;�|��s�4r�ʒ�e�����E���|�L��3%�D?�2mB
}g\O���Zoj� ~6����>���ab0>��qk�j�vJa���Ϋ'XU���=�)Wgu��NE@)E�8�B����B	<���#�s+��Q6{���N|�,��I:E�m�{�{8JR)gp��kYـ�C�!����)�������?��6I����d�>R^*Χ��y��y}�����%���-�������B%:��ibte82���0x���_-;���ff��{����jJ|��t�޴�S�Q/G�$^���T�o�%��e�#!�8N����?�飗_Ek�?r��M�\0�����(���ɖ��jJ�;�Ao�i��z��K�L�x�{���頥�-xtA�E�G][p,���kVH�l�hEP�N��J��iH' \��S�x�@���>ݩ�lm��R�#x��y;n�������W8?8nB��e�x��%���)�I�������8pe��k��+_�\S��rDғ-���Ӈ�I�Ł��̋�r�����>V��m$�Y�Q]6�;=8���|�ᠹ�h��8�IT�h�Je�N��-��t}2�z��?����]�q�e6�I�z���������ޢ���H��a���O�Å�@��v�=+f��N�8�@�偠�����"�������u����i.��אY:��� 6���Jˢ\ދDA�P����EO6]�E����G1�`w�,#��$��T��5��=O%��|�n��1v��.�v�j�>���Ţ&w�&��z�r"K�$��7.����-�> ;VB 	�c��WH�����oh�����2�`�����y3r�
��4��X�Y5q/T`��#h��Ý&恥Fc����_� v�'�ʤ��/���#d2�Զ�E{�?�����h�*�Z{��.u�GR��n5�$ϕH�\�*�}Rқ5�k�t|[����q<GT�nzp$�ꬿ�X{x)�
�%�~����	]�`8
�����舘#@� 3r�š���ڿ(��ݍ�(���_O��4�2f,⟣���<q��
kz�ߕ��!�1�#��)Ζ��M+Z�����G�)�Σ}��'��+���v����j���gA�5�j�iX��b�_��q�y���6Uo�%|Z�緜6nT�z}�n��+5�Y�P+t��@V���vXS�������� ��#��"�"D��kZl��B��x��e7�I6�
=�6I�n�i}\�]��iAW���<�1{�IEͳ;5иwTߘv+*�UZux�J�A��}�*١�$��ޟ�޷o�Q����)�6��p#ֻV�#θ�-��� �;,�A�I3Fxد�Qw�$�,�'j�r'����hVWQQF��+by�o9c�9�D�}�_ ׶�x��N*�M���]�J����ɦ�}�y~/@����?�-�8��B������r�>_W�qyf��^�0w�!���"��A�>*��R8ߘ��7�=v���O���X��#K�~�.*m߶D�ˀW�x7�ab�[��U�UFRC������"xR/&q�ҷ��[?lX�ũ���[��=��b�,vPbC���r��e��c�p/�@�z������Ԇ��H6�Km�x��|y;�J���mm&'��2v\R�ec�]�[,C�1D��n�[	M8��X#Y�,7��`����/�2�)ʥQH���Μ'8]�Ő�h����P�M?�d�q����{�f/�=�)C��LJ��*�.���F0�t�������-1���~6�������|�>�+�>��{N�Ս<�����a���s��J*(͝	��ugxcEi���`��R��%O����'��7�&~����R�aQ�NW���l�;[����S������Cf�B�A���]�#����:��Ĵ688j��p  ���Lg��������I{���.��.�$N�����^	|U��j,�N��қ�s~� ��{�~u�ae��O�SS3���:��J��!�����{r.��d�U���h�_��BZ�A���Z{��k�q�N�3�ڷc��[T�?E�ȍL�?�~�֯���:J2�<�Ӷ�HԳ���=w���i�ɯ�3Tџγ��X��j�������jɁ��Z�7M��O�պ'�,4�UQy���&�>�����PW$Lx�X����?��O~��rN>����>K�)�* �Wct4�h�"�^����O�F5� �a���Fm�y���Ưu߹��St��]��!oRP@>��:��ŧi���I~�)�52�6�|��g�Ir��A��0J[Q%5�O�	�vA �D�'&	�B��ݟ�} ,ژB���\`b������\b���mFtp�S"rA���j�~�kk����3W����S�g����]0)@�x��uI�	aw�C��(n5�>�?��~���O�
��r1����I9;����p
�B��V�����&��o6X�I�,�K6��'H���J�$<��%�#q_�Pq=	/!̮��?�GV̀��Δ�{�k�w��q�LY�V��)*�����ziǐ��l`��&@�}6��_�vI�J��1;���/h	k�g*p�>Q'��FR�K�b��w��[��~YM*�տiDȾ�$Ȝ�^WA�@�>�=��D�o�Cۀ����Ǉ�>#`�Q4H�h/U�r���z����h�v�G��(ۦ"O�Y�}G9Է�?w����eDx�o��v��~|[�ƐD��T�M��9�U� �\S�k(3�h�O����/�&�p4��(�J���r3oYz倓�x��m�X��ӡ�w��E��m;F��Eh��?��\&j�4���D1���\�~q�
򂎘�d�^D*6|�ׄ�T��C����[�.u`v�v2=;��m?���P��Y/�q8��~���<-���^�����J�!�b�u!A%�'�顉�`fsf5�ڌ�t��g��h�\�����_����g[#" ~ֳ�&t��I�#��֝X޳
�ڙ�!-�
e�Cv�p,��Y��CH�ٰV��^
^r�}��8<�%�R)7DG%j�I�>@�����*�_��mJ�%ӣ�y��>�s����p�8E8�ퟓ��&ȗ��8�VkR#�bࡻ/H��laZ?�W�*���8Xa��#s��f�'���������Hn������-y��y�1���� �J��^�Ź�A�)�9�)͑yҐk���������T?"�X���ǐ�z .�NB��1��x�`�(~m�I���1hԡo�A<��K�v�#R5������Q�8�?�0vz��椪�5H�*
$�ϧ0L1Z#��g�<4�/�;33�N2��!�jOm
�\�if]�U�w~u6V�Vұ�K���Qe0ɬ���q�%�H�%.S;�@�$*$j��/�HԱL��8��2��<���̢��k�W�U�j�:9Zpu%�����ӌr�mB�耦x���(�5ux����U��-S��P-��������;����r���a����-&�������G�Ts����>*ht������0U�ӛ��A~#�1�P�b��+1��{\"Z Y{��v	�
�f�8*o�߲-�S*�d~a��7�C��<+1KZ�����Hm�TCw�CCa��wB�Z_h?Є��rd m<7yE9��[�?�X���g-�1���`M�n�4��_�m1,8y�����i���T?W��=A�ZJ�v���Jw�֨:mFL�%{�\,�NC	wbtB�Rv�;Ŗ`rmx{��jR�I�O���k96v<}Ƽ��,�^�B�=n�ǥ0"%[���صO��3Z��Nվ��K�)�c�u�N�P�}��`��R�(��<���{|.�;J��ʻj�#I��'�EQǅ- j%�^�I�B���o�� ��\�e��5|eӾS�d`G`��>�Ŋt��l��j���
p~!NTf�TqZ���� ��q%�N=(C�u����Y�k+c�M�Ƅ-I�a�����G�<���g����fЇl��M/��gJ"mE.�U��$�i�\�Jyp���iJo��P�h�z��g��u;P!�r�tnB^^4��u����K�U��B�x��ت�F�nʖ�C�@�Ub��|���Eo����t������z+-�]]#:1�ƞk8@������!�m�,>��A���1؝H_$ڥ��k�p�^����Hų�r.��#O�PXy�s8=�0��=�l���9�n�^�du���31P�0��Kq� ���hC�[���[���ӱ��y'�1"+,��K��)o
�<�g3V@�D�٣�mY�E<�>+��O���s��l "��[��~0����(�rJ�'�v�ߊN1�u�����A�q��]�r��)=����Z,���D"�,g�L�c�)K�B�H%�r�hz4�[�Uׂ|�;�r�^���v>/����[m�X8e%�^���ڊno����O����XZ��I!�K5T^�ȣ�!ǃk7���
�i�j<������:yY�ȣsd��P�U�}^�Ȭj@��5U�t�:�ލޢ��\�w���(Y�G�u֛&�A��A���#C0qZ7�E�ʂ���̰�!����4d!F�9Sp_�G��p�i�&U�p�R@�+O\%"{�r�����
銛|U���gjF���tuΎ-� zq�$�'T�j��Ihl���eVB'�]tSA%<V�M�^6t`E�}�N&)�{r�.&��37�-4$(�>���� ����Q[P�z�Y��wK��m�sgtuu9�w���:#�m��~�@Q'�T��!�
+�V��fqs��^vR�\^K���8�%��5��gJ�ǘ���slx\/�-���[��jKb�������w�;���ͮ}E@v
/����sÃgU ���3:�i�0���*�UY"�/�������?S�V�ވq��.ɷg�0Xywv��b�߸��1
r1:�pC���O�)PQ;��y6u� ���kC���G���	?�5�����(fcM=}T�O�g�1b��n+��@�1�6ϗg3�n5[
R���������5�~�YGf-���xn��y����3��/�~{?)�6(,��(4��e���IAI����DE��}X̏�*�0���J�+�����>�C��`�ޡ%X�gއY{�<qL���Z+�����>����#��^�'�;��!�CYK���GzЪ'�,�{XO�T��m��� ��&�gvVI(_9W��Ҍ�w�#�Kp�'��9�#2�V����G(�¸����s��H�z�.%�Fݖl;�}�+!�EO�JɕX~��e�L*�ʾ��vc���i�x�1ѥc��-'a�E'�ۤ��'N-/��d��E��p����fK�hױB���>p6R���l�=i����\\u�������,�g���ՙ<�W��Jx��`U��#�(wQ��ǿ��ѷ_��1��4����}P�&~�th�(�S�(���hWz���\������85����|:Rك�1��321���f/IU��dI�~%s����19��b9��L�yLv0�An��.�2��ɏ�X&̓]�iFXA�ݬk��u
s�Đݣ�qZ�`h#W��,,-�Yxh���l�Bd%��ع��7S���x;�b|ֵ��_���Í�z��p��;����A�E	��o)OB���2�7o�ߟ-�VC�	B(����G����$Ϸ��^K�*)FQٳ|�ҥJ>�$2���ݱH1<
#v��,�.k�F�}�9g�Zj_A��ιu|o@�A$��M��S��h���V��'4�X�	[���V�;,�t���?uơ=µ�L�P��i��0$���\׫�X<�Zb&��ߑ=^[BN�ǆ���@���h��e��3����1�E[���	�����D��tE��z@���D�~��V� ��v��8���@�R���Q\���f��Wۅ'dO#�[#^�z�(44O�G�~˄m�Ϫ�J� ǂ���J����K�g6�jg�33��#��C[ݎo�ʰXY�c(nB�q�q�f�N3v�bh5)�LR@lQb ����v;!4	��ϥKHeX> ¬�'�}~��=��q;�K�ȝ���NλFV�)-����D��^Ͼ�u��N�[$6u���AA	��X_��l�4�]]	=�
��a�F���%���1N!��*��:Z�����-P���^P0|H��^�Ǉi��)��k�-4���P��k�n��ʽ�Y�""[w��x�rU�3Ԛ>L��jK2RT�2[��\k�����Z�ˈ�D�[M�u~8Ìh��ooq9oCN�*#��P�3@�b�|F��Yi�k��H�43H0�4(��a�)����,�.�%?@�Wh>K�8��E���>J'Sc�=R����BO�j-�כ���u\�{��8�ZM]f�����
P�A��}���W
�����^���3F,~��V�����B�0�!|�E�M�M>C�i������9F����:����X�\N�9����q��C�>�rm�]v����,	�yu�m��!�e��G��G8Oqy�S+��c�h�`tr����&�-�tSҦ"�r���������9�)���9&;3bF�u�o�A���"��֠���-�]�&�%�s������Ì�w!t�v[.��H=�u�ٺa��A��P3�I4D����Ѕ`��������^Q`�g,x��T��w���g�
xN�޶Ȉ�~�LT���4U����[�ș����� �#�4h7ˤ]F��m����O��	)��~���(X8�o��z7C��`8G��q��ʦ����6a�9,XJ>�a�0�g�rf���Ih���f��Y��5m�l�G�o���z�YBqP�W-����HhK�	���f��i4
��h�w��:�_\W|������إPMSm�2����?��Ku�|��^���l,PNɰ�Xћ/&�sQ%� ��_6S����IE�`ej `!WUw�U����ȴ�n|���F,�2�0����%Bڤ�'�+�!����7���2ȵ�Et��#'E-����i�-���*��A����[νq�𠝌(z��X�`�|����2�.�z��6zFж�����*#�I\z�~Q���������R������y����n]6�;c`õ�h���*�����>���I3�}��n��"w`��q�����2`�JF!�f�Z�3�-i:�1f������ޏy�4�%+�ж���j�ܒs�����P�Q�J��P.�B<MQg���6��&��Уg��S2�3��_�� {�����q���@<ɘ{G#���r�����>'���θ4��ȮOm�k2��V�؀�#~�jW��:���&0�L�Ja�y� ^4l��P�]�Kq�O�ǻA��⮣�i#+J�ͪ�W:� ��^�\����zߒ3
���&sd�=�*��D���{�LG���S��]�1;�r�>6J����)I����(W݀@����G&��5�)}-�E$WA��U_֨^$8E+�ETs����j6ڑqTE_��Iy�'�\�%�ͦ��F%ա��?5�S�P%kowiD��8���I�wnb+ǖ���?���Y�+����G�H+�.Dw�8@�?�O�/�TYK��lS|�n������FPc��ۏ�lìR�:������N����nxj`��rPC *�GR�&������_�1�&��E����&������'�U�5a;��\f�~��VZwP�q�r�ڑ�{}�	&Uz
��\Pw[K���)ʓ���^b5J?#�No� a�v.>���U���ᖀ��4L4��P�2��vbO�w�����r�(:@MѶ<��-2s�E|�pՅ۰F����3�F#���.����RD�T%XNO�<���$ʕ�3�H�se��I�<��>CO��&���Vo����A&����Mll�Ei(�a_��S���� 5�UR�(t���<ڝ����@i|��)����&�n��V_�����s���sM3CkB̜>�A�E�>�|�N�?��@'�g�����r�P�F�	\��y!4S�#��xK[�6�A[?��,pIA=yB�#Y��q��s?�D�ְ�Oe�w�E��9�m���1D���޼����n]�FRj����b�@pQ��ͻ2�D�=}AI0��(�e�,��[��o��C��� S|�-V���
A���(�
��,QI2�)[f�1j��+m�$cW�VS!�]³.8���y4n��9�t�i�y:v-���v��i
���8�ѬT�U&C�W��Z5�!����`�v�kmԆ7bI`!G�H����yK*��o$�©�㜎�hV]�rXD��;m����w?�E��cW�Uu�o��� ��U�ì�}��!QV8Q�1g��d:�ު3���DY��+�ΰ�t�!k��nު����"?����Z����AK�ͺZ�Q�O �>�@�/Oh��P�asK�sٌo/f�C�x���(h�:a��8��,�	�|DF<��K�/"�d�6��s��".y�J��։F���Sb��	>�����}���HA��B��;�s?1��#m=I��������,؄Sל����qV�0^����N��P 5h� x�Y�nv�d�ʡk~d�,�m���f�S���q:�<)�l�z���diR�[��H�a$��)d���.�
9Vz���8�Ò P��7y�������
�iN�\Ǡ'�촚2s��Z}��-g]6W�2���C�j)e?cwo����,�����-"��i0w.� dXA���ͨ�� @>'b�j����U�M 
�N</I�f.1w�L�\�Jr�_t��۩�*�*Y�U��6��|F��@�ՆC�]@}֥��z��c��X�قM���Q�H=��Ϲ���AT씑`z}�&B��D�T�ӽJ�ƌ�N�TI�d��6��S�3$��[�v��n�:4C*fD�/nC�Jŝb�,��&�w?Y�����Ӑ^n;��a��~��=Y����=n���|��\ѕ��M�Uί��Ä.v��G͑2Y����+�+e�����smT�(p�.��y؞��i�a�) IA؊ɢ�i�b2yR�k�^_f<��'D���*���	%���@[����zo7l��mȃ�;��kō<�.\�Ԉy[{��@j�_q����z��|��K=fd�Klw���t�_��E!?�x�S
84��WZ��>�DЎ�6� ����k��E���;�,����~X�1p�VX$+��jN�4	>z,B"݄#@?*0���$s�8�笿j��
g�|��y���=������U�����f.Rp�亳�T��u�S�k�k�����Q[_b��{�:[7_?=��/�QG��цi�C��\�J#�T;9��@][��΍�/#���T�6ּ�P���S���o�՟���1��q�fOh-��h١��D`����E�߃-����7&<_:�+�K�C	v�J�8�SܞK�UiV'�fr���ȶ���)��V�cb?h�i�]g��/�C���Ѥ��z��BF^�ٸ}Q�������EqQ��44-��Ѽc�=6�L�	F�ȓ/��Z5hޓUC�u	��^%��'oBӐb�M5gop[+9�Id�`��C<�Ah�\ؾ%�"r�� H�J=C*�#*��H�E�����=�>C���]�?

�T�|���Cdl@���9PT�r^�F��J�b�5���jt��/'n}Z����]\�Bx�󿯲�~��6�����g�	*�['��ė�E�v�b�	x���w㵭F�ͱ1�Zqr�VT���n���x��D��-�M�;�$��u�K����W_-#�UB��~��0w�|ȅ?�H3d,�������.�%k����Pi�Pi���˽���(��,4��}�h�1����W����w�� �r��Ks�e~b&�oB[�ŵ_�����x���m��@�j;Y�����و4HB��*)�4��:�˂�j ĵu��9�ME��\~j�R���u���|f���$;S�2૜��[��z�ޯ;��a�u��O�T�|�2�)Ku�tU���R"Ǒq"�I�a�K����$�8��w=��J+%�ذi�	��,mR����K��G�ߑ�,�R�v{�_�qI"�0��>I
�sb�[���g���F���z��yV��%�����砭}-ЍI��F��f|��������F�(_�H?*s G:��ɝ�c�ƇP4HQj�N�~j�풲�}n���?C|�|A�qfC�����0:I:y� ����z?G�vxI'o���6��f���y&�k3{8di�� X�t��8�+)��8�C�ڽ]�9>�9Q�2�����ItӜh�n���N_x������2�n����Խ�B3Q���8�r[D��}���P��TN[NHp
(�Q�����;4qyG�H�h]b�1�j�۪�k�V�x� ū���2u3h��E1�Nh����{���76f&��JI� �wdlk����w��(�-Ш&�'-"�>�͟��bR7�{\�� 7�Q���J|b(��%�Bړ}c(+��Z�K�`�c��}b<F����_{��0����m5��̥�~'�x�m�[�a�(���R�6	�ߺ&]��a�a$썅܌�����c��v�Ӧ~4�{4�ج�O0��X�r��r�Zv������� ���X�z����B,&T�(wR��3��"��/u�|� �+1#���ٙS�s,	�$��z�u���Ɔ3��.I	�8��wzٿ�	��z�;*4�x�z��jy�g�U���N�	�����)�p�h�{E33�"",�E����eN�3�fl��U�-�+���[���Vr,��m%�d��Uz��zkd���_3�D2�@�!���Ꮉ��%�pF�~I?&���"lR���h�;�����C�Y�=Q����/��6����Z>�*�����S�I�r�.P�"ߑ>�wI#I^��63����9�t��ɱ��)̎j�>}C��w_�
��j��{�H�<�$��)$H#���U"ki|�+���KE���z�|���n>����!p�Id���PT
�uo�)�0�����a�h͔����gW�ۇ֝�En-�EB�H���,S��<��eV�BK�@r�%��w�3�T��J�=pm��:;��B�a��w������@A]�iL�T���c'Z�v *j��j3�y�g��'�8z ��z��(�?l~.�꒘��U@ZZ��'2C�OQa�W]UN�C��F�0�[��5���7�y�Wt���0�5��Y��RUK���ȥ�1]�͋V��ʇ6ۛ�lߝ��]f��ϧ`P̜�ۊ=e��[��B��ݎ:K=׵�`?\1��g~���{���
"yS8V���#���y]�TE�G���.�%u�����2W0C6����:1H��kr^�KϏ��U����Ru�i�'|�1y�g�ۼ��{g��i�Т�B��s���V���2ԃؗZ3�㏠�4�f���"-b�P��▍�ReY��G$�/�Y|����S���lR��_�IbW(�2RnI�\���s�=~�JDG�'��9�b�L*�]��?����cy5�b�_��m��l6!_��.�����U4/�T4�`$W
��C�sd8�~k@5z�J`X�����98���L��Y�0��Rq�Q:��9|v��D�{���S�0��癧����LzE5Jݜ�y]�@S�G��t逥>��֗�Lf3(ܯd���I~w)a�h�ܥ;f�Aʠ�r�\�0����\�u����e�\O�;,��1����"��}�,����V�#����ρ�'�ˍ�k+����e�� ��uW���5�|�;��x~b�!�t�*z#>�����ʁ��}�옏0�|AW��Ѝ)�i���)�$8�b$�Ad�}�`�NC^�NɥB�g�kM������G[=�Q g�~�9��8��۵f��qf�2�Mo�joqX�a
�����F��)�]
��K�Gʐ��5��^�D�ŋ�j�3�Mw��F�J5�Fґl�R�����Nu�a��#���!�G8�+J��X�M9��L\ϒ�fIvOE�����g���^}d��Z�C�\6�.S��	z$����J���0(_l��_�>o�!L\O�P<�d!��?>R^ec)�_�8v�	6���W��i��#��Qx�SB��0�R?)�:o�N�9������j�A�	%��*��!AS@T���8Eز�J�XG�����p���: �u�.;�6|F'zm�ݡ�Mv֗R�k�~���9�,U{�o���ƈ)���E�4q�HV���W�|8��N�_GA~��,�a_f޴�x�4~���H����w٪��#g�y
�N�p1�m�2��q��Ya0�$ ;p�˳�Z�F(�f������9F�H�ʒ,Q���*j�y���9$u�����Wm��>���Ͳb8,�$�n��Ą����yn�^}P�w���a�ɽ�p���:u����L�%�q�V�!#Yt�2� �`����}�}���W��»�{��	�I�����0lv�X���[k�m��z�[q���{�ˀ>�,G��I�:�q�hm*S��;����k����R�k<E��X �!�{>�����_�ͭ�[d���S!��b	yU����i�s#
5T󝑝^��ˤ�3�3Q=8i�������	��`�y<+�|.���}����^gɅ�Px�ƭ����P"�q���E�K�M��Y�
�H���3��R�1�q6���:&̽BnLU�_�WR.㊒��a&������vF�.K��!�B���z|�|�,ԇ��F�^]_s�N��B��r�E���]77r��2P���Y�k��U��V��X<h�Ir���,Z���t�"T�yN8(�1B����/��Y  �ޞ;�(��EG�Cc�l �Y`6�w�K�#����y��.��ƪH��^����X?)�};NC��Ěr5@-�%<��W����l�����}�O���=0m�u�g2^�?�{%�#D�)�1�{y�fa�i�T#�EA/�%'0�^�[�B\��P�u�mpY��3jұ/{�ŉ_�*j/&v�9���校�k�k�f,W7As�;�Թ�g۴���F�W����Ȉ�-ѯR�H�:No�V�1xD�w[��Y_�f��漉��R��Jk��ss��N#�&�Zէ��x±����̗��Э�#�=���
?��P���"H��z[�\�+����+e��˹��|@�J�yT��ﮂ�1�[�V�Z�	���:�>���}���v��W��5��޻n�{0���2��xa=i[Q�����~���?+>��x�����<�{Fߟ���?د�f���'cE%�*�{<fth�(t�u1�죊�u�%�^D�C��Zh��yC�gw��6�l)J���|��o�xn����:J���ȯ��jŇ�|��/��.�����%K�t�Z��F�WyԓY~���r)��NVQy���''9���'�~Ec�a����,��U�n	��* �Ev��6�U	��Է*���}�~8��g���7p�-��ϴǋ��~x*T3
�76m�lMɸ�7ց��b�@8��:-�v�zQ��g�@��/��צYݷh���Y/U(��Q��E6ɹwx?�I��7 �Tpy�:����^��_�\S�w��`������S�
p|g���6
*�~������t�1w~g|��(��l%Ě�XI�<�M�r7���+�Cmz-b�jN��_�ՠ.�����د�"^�}���8�	�9���s\v �:��4h��$����.Y6L�iY������3��*-�E��A͌�/�ɐ�N�58��<�Ǻ7�W������[K=0I���6"9ø�U�j/G��uʡ!ȥ��%T䀇��ϊ��'F����޷"��z⒊�[��j7�b�oml!籺�z�j�E�wSwk�ȭϙC뫫��`םR�M�Z��v0�ۡr�w�~�ӻK�1����O�pq�Y�+��
ǁޤȝJ�b-LՕ���<z�K^���S�6~�4J�c�:��+� &�	3����+,>��8#%�J�-�z�tfBW2��^%��ZoB�zŏ6e�[�c:ǋ�AB�#r!�6up���n+��j�y��_�QR��x�I�cY��g�yͭ�`82DP/�����<��ɀ'V,y�,P���o���^�����*%_Њ/�)�9o�r��Q�CsdZw�F#�Aㅴ?�Y���w�+����z\�V+�c�J�H�/��K�5�����k_�<�{�_д�sj���A�%��V>��c�Xv%h� �sQ � Y@�O���OFq��p!�Ⱦ��	ƻ+�J��p�U�gJS-Y ���'�5�gKm��WuEU�!�WQ�TԹ]��l�t�~�
�D����z��tf���r5:�k�`�1�s���� ө41�{�[���RI��������rnW�Ѓ�h8V��a6P�MtQ<~��D�,�ͤQ8�Gj��]�*����=1u����45z�f��&D�_}�s���~���|�Ĳ��8H����P�lK��_��П�@}���?+I��M!��m� [I~�T�R��X*�He48wEm&��*�oғ�!�2a$��ë;��$�4P��m��\/�[@� ;��?���EN���xO�S�v�I�jD���=�E`c��(Qx�F�~^LF�
	�j��t7����E�I��h���s��Y��5�i��ܟ�;�y�k3 L�����NW�vBCm��4�9,<��AG�������^ǅn�����rhe����0�=@ϔ:��� AF���xQ�)��,�N���[3E<,`TƵ.�&�.���ƛ2�4@8n謓0?ku!@�2�~ߎ9M���́��;�#G��0�^��c�ϻ��i�t{עD$h���r*m��6���<Myӱ���%������!lF��ņ��`"�� s�t��n�H~�DhP�0¡Ck]v.i��r���m�~1bc�U���7�E�8�`�%������ѷ���w��DK��X.�4]����$ع�Lf?T��z�2�gN�ލ�M����՟��VR��s[��L�C�+�����Ӂ�5s1
z�����3���nG_G>�v���wi�zn����ᡁ��e�O��<��@�ɺ��an��>�����pn�fU��:8ñE �/-sب��R�<r��,�?1����a�'�&7f�?����Zy6iW3��@�mJ�C��2�3��gZ�B��m #�"�ћf�&熥 ;��(��	������|�1EyNeV�`�||�r#_I@3h�4�(L�Q���kZ�&n|��S#�{�����O\1���]��o�P����у���)H�'�� �+9����W4�nuf@>�4xAH1-ɡV��Q�|���N��ji��a�F���\i���^v��y1�	�ۈpҌ*C��۱n
ƫ�H.7l��Z���3�(�-�E�dW��i�l�V���������:���<4�C��3���q��D/sM��pu�oX�_��c�W��&��v�,M�&���S�����w�'��.�b9]M���i�-eи����a�}	�u-��n�O�~GK��\�B��� �B)&Ky[�e62��J��sɂ�p���ح�7�Қ=��v�}Tj�����	�H���;��M%� -�l��|<�S�%~�Ժa��ɕ�WI�y����#:<<����MP�m	t��=ʱO޵'�`��n�i5�ء��>%�xO����L���%3�|%uZb0;YKEi췱5.�H.����w��ݲ^�>�J�j����N�bS�NF՟a@���� ͌���F�_�E���'��j��x�h:!��=�~׺������Z/`��"�D�o��ՠ7�!]L#�9!7������ڔM)�k�*�HG�iC�솾��V���؋��<n��*�R����Mᲅ��IAڄ��O}�w_Z��s7�M�h��r�W8�#a��rd0�%�C���ȗT'��,�p,+<�7�~��p�њ�6Aճ����i�
�E�S��Ā~�[k���Ʒ��b�|���*A����uǐ�"��#k���㻨�*��:v�Æ6'�.!�7dp�%ָ�{�3�i,q�m�_����M��s�O��/Q��ڲX"U&��j�>��[Q81�4Iq��s�t��t-�^����^Bj9�g��y�N���A�l)��]b`��&Z�wym��Xg��J�$Q��z��gF�r�TM����@ ����Q� ��A(�`>�
Z��b!���r0>��1���-QvF�����Z�/�G���D�J�|�\m�2�P v)�I������nó̮R��6(Ծ>�cE�p����6zO�PϚ�������iダ��}q��pq|��������Ll����Þ� �%��(U�gd���o���`�Ŝv�pA�R�2����qC�q.�6m�}>�Nj�!���1�P��rv�sٻ�C��k���9B�rsL�b|	�k���K�O[������Ȋ��9�Üw;jY,��^��ئq���-�M�i�bL���)�O���!F�H0�{��}�X�Z��7T���9`1�Gr����Mt��ae7?)���WN�s�e�F �{ѱu�st@�H���	P=���P'�F�[��_lc������q��}���_��WĂ45�7�}��\����@eLȽ����3d����g�a}q-�
���m��H���7�K�Yq���
��� ��L@��J�_�$^��'D1�
a�jm����'#d˭��M���3�a��q8�=�x��9�5M͉�׈VY��5c�ݤ4�6ݳz��rЊ�g��	}�%�ú���#M�Kb�?2�f��!��Ĉ����|MT��.j���bm�jw7�Egc7�г�#c�_��J8��3p��al˂!����- ����eX>�t��YC�]6�#[�XQ��o��}%ƕ����Ƈ!a:'��780�n�mˣ�CO��;���d�� ;@�i��)�*�xA��n�`�H�i�-K(�"�� ��780�o��6��T�ق��M�b�	�ψP��U%��Iv�H)�[���\�{�g~�Ծ������ Y�M�颱��v�{�#4	���Lo@��6�?��ABi>�0�=���L��8G��
{���1~#���*��3	����](�T!��\L��͟��/��r���Y�(oeg�ӺL'fd��t��f[] X!�_�J�x�q�q���|�֟ο�m$�!��wX	|}��eO���]�MO�C�N�w'`�l3���%���ެփwb�]���� d8P?>֑=oo�T 5�Eи�K>Y\au����L���j��]F�~�����,��r����1w���q��^}�'WI��d�L�us$)T�b���AV�^�1Y��`���R�������y]���Qdoh�m��:�3w������4����] jDK~�k���슊I>�,
�'�fF����	a3�&����,)�����<tD:�!V�Fː ֝/Y��Z:��.��aD��U�4.�r���ѭ����"OC�^U�&��8�_�7�^Zik�Nt�ş8=<f*�+�,4�6�#¸p4<��e��t.�5�x�\L�l�KB�n��?Ԗ>q
�+|�;����P�k������y�n�vJ��^��)QG]���I�ԦB���̶��u��	���eׯB�Wu��	q�撀�6�������b��Ұa�J���D�Jp,�Y�o��PY�������0�m.��3X-jp�
D�~�y��b��?x�.�����;[�Ԣ	I���c��_zX��dT[nN�e����K���~d�x%g��-�ixj1�I�����N�D9湴� � kT{�L�\�ϕ���tq�{_�Q�\��������E�pQ���jXeI�euc|��&7d2�Sx���w�r�?:E;��.��'6�r�����}��U���Ss>�~�Oa�z���یR��0�OɌ�w���fi��8�H��;�%y(��b�^�M�]��ƨ��2⩬{�_��hvq�o�;�+8�QD�
���^N`����������.$��a
%Im��y�3��k?ji
[�\b�V�����}�6�q�A�e�9Ǝ�8c�V�_�6��LP���qk�Jb��_�9//�'�	Ģ�ϵ���WbGg^y��ˡ�X��x�q��D�3Z�Bӷ]�Jv����>�����fQt� g�tEteW!��X�1h�E"��A+`��g�c�AE���l���x�ECe�G`P7�!<�r��%�Ǵ>�Vc���I����f�#�?r'���ߗ�:U���c�dA�BJ�X��΂zfNB�z1hb]���4vJMd2+q�6�k9��]���O��&���Wx6)%u�09m@'�>f����BPZ�_z_�1��a�4=��,�DBAs6���.�A5p�Ƭ�6�a`�z�[m�LhS&%�f�� eZ��b1�
���?��2�*��[��){8��sJ����ف�nr��ۻ��j�S?7*�t��|�?�y����6y��/��O�B�A���[��t��/O�ĥ��PX�����FQ�(J�R�/J��|Z��I����Av<��ij%0 �"m>��+o �����*�L��fCD2@�k�w���S��^!U��6��
]�ƞ�ݝ&�+K� ��I&)�H��7 �7ͷ��[;q�����j�v�'���1q�eB^�t���T���3�c��Q}=VE�i�L�!���i`���)�r0���C�O�{���5	J>�ur &�(��KH��2m�{�4��4g�}�A'����9	���\��>J����`7�U�x�=���]D����=Y-ڡ�|'���§ؔ����뱕�Qղ���P�����m�5�?�3=3s��+�I�);zA��e�<�Q�b�^)�`�8D=Y"ftz���U��7�č�]p�ùt��H�>7 f��B����i�}Z\���J������ka��zA	�8A�<!}�S;«��|zM��D�cRE�)���(鞨_kK�L��B�/I�oˇ�'�bg���e�AN:X��4�uX�zXi��C� �'�g�g�����ӈ�߄l�.��:���,�@��AgW��Zk����g���3�� ZQeھCW�Ƞ^_����Á������ӽU�H	�y@kd[(v,�4,yLO����3�YyϤCF%J0
�������yP(�n?}�}2�G���X2��_���p��Q������~�gj��0��v���|��"�q��T j���QOɯ��/���b��*��ںV<C��fV���G3_ G�BCn3(�ix�R)
H<���u�l��Qڏb�W`�P��Qh����`k� �d�{@�bf�P���k:����+YފB�8*	9���d_4e��W�:nÕ�W~�2T��Mi��i��_� l ���JÄʷ�v��읃-��Ԓ�a�j�C��:���D�$s7�(A��N������'��N��GD�Δ��{}8�XfЭ~eR��#����ݻ�w�˕U�5�zfy@R��G,��G<GM����"����sdI؃]z��bm���ʲ`��-Mߑ1Fc�/�qJ˿x(w�l�`ܾ���c�N��KB�M�[�"���J��H3��M.>���w7m���Y�>knQ��O����2=� �
0����[�j�U�햋ի�X��K!�?W�H�U+M���->=�.�����|٩8]$��v,�o��n����QX:P"�+Ј2PEӧ��&���TMr����c豶�(tP�Kl:�7hq5X���l �6�����0zGC��N�6.��;�c��ey�g��[�߼=ݻ����`��w���k�Z�WGy	9����zK��Z��CD�g�8i9�1"`�fdO�v����Y�Pp��H��4�_D8T�_����J�J#��(�&����V`�~��' �,'"l���9�5�0���|"�z�É���K�)vp6h���b�Şz��܎+��,� Սg��~,�%C*�k���v��~���:����%H�}JT�<���� �F\T�+e��!T�V���|r��+ִ�r��i�WD
&�c ��GG/7Q����f��
�V���"~�����͌�j���!;�Ix�ԧb�+I�e�����:8���"Σ[YIX)�Ƚ4���u�IW�����B���1�ϳ��4�W�nH�{X��)B�ƈ>yn��B�]`�e�}#���ڞ�pq�[���̣�%����v;����j�q���['������ �yu�
��f�s�Fj�^�o��9zx���U,#��=���byƆ�p6�LU�Ns���Bo�O("��0��'�U,'P'ԣ�qd�_�aj|�n��IE�eav�@������������ë�ɕu�s~m��<L(�cS#��d&TfJ.�E���F�k(inx=�;�fJ�C�Qjwk�dd��t=�B-���>Ƒ���2�����2�+�MHX��eE�0����h����*
�F���2cry2w��۰0L��]ٙOYc��n�=sr�<M��,����N<bS��r���l­r3Aߺ���|�č�T��I��pw+��kK1t�5��#�XI�Wc�G��`��K�\gh�h+f�4&����"�U�mP9L�dŌ��c�X����\���iK��eBd��������L~�:Zye���c.`��*�ݚ9�o�O���t��`)�w�c��}���\Hq���]��*��*��>�m�/f�����<瑅	�.�p�u�"!����; t�a�}@�d�z�t�Q�.�Xu?�)[���Ү��35�w�jCﺬbP��	�o�A�i�i�H���_F	9Ʊ�8�'%#A ��) fj�
��n
��Q��\��������A觛�47W�kr�H��nڋYĶd8]c�����n5��-��z䃝�	�W?6
�J|!F��J f ��K΃����
?,�Ʀ��!�ŗ�3�� ���w�.P�'���͓X}�M�C�H�V�,�f����LȢZ�qRW"�u������B��-�,5�2��uA�n���{䔉����la&
��jij����w�,���6BihG`3Q(�Lא�pAz��==�������c�b��%R��:���S�b䬘�_� �����n�T�����j	����4�$Ԍ���Mi8A��ޜ�$�l��@�>SQ���	�y0���n_x�_�P���J��E�⪑�j!w�"�����ر�R�Y�ɍ�>!�"���e��t�Dp軘я���&��<��:��`����������!�W�ʐ��O� ���i7؇���t��i@�_l@$y�4o�el.h^�<��\!��3�T��J���dVu�t���b;��&!��2��Xb��k
�����������{i��(�Ҏ��%0?m/��r���h?���@��_F��ԫU;�
��:�*_β�]`��^3�a�B�;>>b�3��DV��b��}Mk�8���Ų��k��%r1��ropn���P�lk����h�^�c�꿾���D�aL�Z�Jmb(gy��x����av�6�U���x���ͫŝD*=�E;�8K-��bq)/a\K1_�2������@���^��$��ҁ3��e��u��A�1R���x%D�R`4%��+��<��Ep7�Е@��Z�׷�R��R���եg�`���l���CnNFX����~��D��=��7�E��ޔ���XH�~��r���}$3�k^���̌;ʈ�y�%���5%�h��W��H�����Ĺm�7�����G��;N��n	���:ӉK��!d��dG��#AՁz���܎9%!�� ��!SU�M�>�I�����UZ.��o�#Q}Oc=I���<H��"���D`)�;z��M�\�kĺi������wMFZ~�Ԡ،�y:�)I��D3d��s�.�w�Ec�M��o����6�1FH�1�2�PF�U���d��:s/I bD�j�Y��)�aK�y΅+�&��?vZuw�� ;��n��㻐�%�?���? d�+i%P����J��+=���J�C�Ͻ���B_��(V���h�*F
����Dt��H�(5����|k�������JIo�Qn�R�*A��z�[>2^r��∟�+,�eө�C���׆���J�Z���U�1J(�ln�i3���4�(��՗��c˞��N��m.�S"\�3PL?�� ���!;�����2*�����wP*G6�	�c��P�F/�q!b�^fM��������C/߽u���APkp��n���B���P��:��A��Dh�ec���	�[ՃZN#��@�E(�]c�*���
/劵���IEr�'���4e��Ӯ�����ݫ��)���gh�ԉDd�*�6tk�8 ��t��e��VY7��'�Li����x:F�V�����]��K}����Ŀ���F�Xz�­��y0� O<�2���5x����N���K��-�����\��\B����m4%*\XaT�Z���+_5���@ ���*���א={��#m��jd2�g��-K����Zj+U���39yΌ��Sri'�%�����Mج{A�����{����λ<iD�O��4I4��/���)�D=+k�޼)����h�x,�l��(��S5��������3�w��=El~Dc��.I�2��L��[au�W�ص����^B�<�re�>�o����P���D��n&� K5e�C@�#��e�`,_���b��Ȍ��[�4f���d�E�e���S
��6O��Z��������쇊���D�:
3W�H��8Y�<��L# 0����+KV��o�㿳�CyO�Q��i*45��Eh\\�)#ŖP?ݜ�c�M�mA�ġ�I),�k�>�D�4lA�:=�aV��=;/�+`Q�Z�}Q��+f6r�_��	��`�[
 x����c�o���e/i�פ��� ���ܚ���������Mk�C��/Oo֪'��Epӏ6ŏ��_k�WPܤ]3�P)'5C��{H?������w*�nk��4�y�P�-�7
�at�
��a�������Q:]]n�gxc^4�S���i ��\Cu��
��V�'A��O��ց�X�` ^ne&@���:F'7����^�@44r��>bc)P4%$C�"��λ��� �T� ��Wm����82u�q�!�[�+A�X���tu?����q�.٬ҕ�\�c`YBN��w|�@t��3�^�3��K)(3�J+E�������γ��+�G��7��W'-� P_#%l �a�S�(q5@=v/V�YdMd�-�N �5Λ�`�E� bA#<��O��UV7��S�b�#]:�,�·Ϣ�+�b��)��ӻx�)p���M��w��}T	���[���̘�9m�K�̃��X�$&�i�_�n������4��nOOn�(��Gv#�ņ�q�����b���Q�C4�k������䵪�Y���Ǫ�@[�\�tx�n����B=Xw��D�>=B�D� �t�҈s���-Z��+;�⧆������ �	�d�/�q{Gp�؏ɻ��+T�P��'눅mmu��Y�/���Q�rB�O :_���3e�:^'С��J�����}P ��y��2�� 9���J�k���L������]rϻ���=�@��2�K��n}j�z��,ܓ��,�)�7�*�o)�!�������0c�@�X�O?~��5O	B���"5��)UGs��t�+D4�vw�3ud�"���\�Ϡ
�?v��)7˜�������ȉX*v�:N��]V0/v����:�ٛy��0d˛P�ۛ�F�i�,V���U�s?2뗏u[�����Ln��^�e�d쐢�:qFk��w��g�sJϑ!6���t!�*X�<l�Iv`i�j;�K��b䪓��N�zŭ�C���&����&*Q�)N/$�c��Ŝ�F���@+p���:�MB�k�[�v&t�O�m�`ޟY�a%�A���4=���s�9"²�?hB�譵̯����9խ�Q��q{P]�/	A�6���Ip�jƈ��������&#5|�5�������t>�7�2L��A^t�Z\�X\�#Q�-�J��ʞ��㎁�%�L��E����<��BG�F�*tu���8� }T�$�R+�L�;�8�� R��%S�u�i����Ln�q�,ɷ�E�@�� ��XU���}��&dxf�C�RK�����Q����ke�g�nmF+�j��6�~������>��nDv lb�i�l�u��F��&hHY(��"�㥳4��:�ˊȷ�l��xp�J��܍eYhUu}I�?�! w5��g�"C�
<�|�~4�.&Led�˧�P~Ź�RE�	��QY1�2�O�¶^jN_=e����~���S���/Z.X��</O�N�4��z}%ð؅GaG1q�>��y�b�����_\֣��-�Q�NgQ�~���\�9�ѹ��Ɛ��]�{N�I	��Tl�o���H��4,��+j�D�-�?9`�b��	HȤ���0��?��a<�9���|�28�>�b۬���f]L�w��1#�z
�2�4�-�#��K*���N��iWb4��u�*���h�����=�x��?$[i��j����v����ZJ1N_�f����_,��۪��u�Q�Ҩ�R*�)����44�Z�M�i�
�Ͻ�ԣ� (ƯdG��zDeR�����yRR��������P|����y�Y�{�05�� �ɜ爻Ar^Qݓ"����V^����$_#�����\	j�j��ي�e-�݅#h���Y��5r�f�b����_����N`B���tu!#��L"A�i-o;�yz�GLy�\{�y�R�p�G����k]�'��|Rw�tlt8��n������D#��+⵰���c"=2�Q���H$jEC� �sڅ#@�-����&��;�P_U��@?���%��HT`��ς}���2Mۦ�͈����È\���'�R�Y��ļ�JR��ك����Q%�i�y�?������o�W��A��B�w��A�o:�˶�4��=���Q/�Q_��~U��/���Mئ�Q�W3)��I�lduN�	� ��fhV�����"x�$,j$i�J�c�#!A���N?/J��5�8]��I9���eR��� @�
�0r��!�QGL:�  �=�����	rbDp�a2�b^@�v����J����MU�q��m*AsEŢ���t�'A��f~e��a�A��}�E�\�S�ë��h��PV��J?ڈ�B�'����h��|9NƝ`0���x�|�j��������"䧀����R
�Y|�o�6q�K�� r�1��/��Dq/2ቘgQ�'WIU�0��,_���'��V��c���W���Lɕ��{�L�V}�n+���=,�Q"�3��$�w��M�\cLd���9����tY�.�\��c���9v�P�N�J�Upn��O����#�u��[�$i��_��k'����7��~�����%�|�Y4�f;�^j.4� �A+��k����4�2cv����J�j����h�p%�;p�: �����_d�d��? ��C
_�eL����_r��NE��S�SV�Й��?�\5� `�[d,�B$�g�̟RhB��Ї^��Q<Ջ3��t�����+�Ik��������cU��������hC��=�U�7��{#>��Ī�x�Ăz�:U=N�L��ܦ�M�A��H��9�	��Y��Y9�<�r_��D�d]6��E�B- vm8l��tJבE>�EP�@v>�<�(�^��ޑW���6��b�W����q��^N�w�9��Q+Q��;J��Q�ճ�\�Gʹ��ͭY��Ȭ��S�U��&>��챬+�F����0�쌊�3c�%�i�>��"����z��3`�F��2co�R�#^��~��	��������m0?����>�����.��u[�Ӡ�p1�s���k�6��/��oL��9��g����Ta��u��tZ��u]���F�y��UO���c��d�*�U�U�BQ��(��[���� �q�4I�9��7�j��i|� UcT����k�5,Ɇ��Rƴ���:���b
,�r����C�͞뚃^*����Fh��X�"��1Y{�x��k�<�3�)�I#aT1�����k�Ce�+�6�(fL\g`��N�c����mUB��z�7��ǃ5Kj5�m���� /@����£����)j��[Fɏ�d���N����7���gXJ�r��������D�6�4oVٝ4N�<ю�^�s�;���s�#���A�0�������c�^/�.�b�j�ܡ&�����&�|)
���Oa��e�3&�'F�h��̘��y(��S/$θGO刅C��xX�g��v�h�y�{W�R�ޘ�7�&U)���B���heÌlӇ�����뜒[���$�	�����Y�V���ڤr�-���}W�C���g\l{Xܮ@S�ف������!��'ʺ�Z�����"xxd��s�{:(tD�$�L����a_HΕj#�W��9.I��'FG�q/?� ZԻ��g�5�с(�u�z��N�W.��]j�8�0���"��bK@lS��*�JL>�T�� � #�
�E���?*�#ǰ�1_| ��ѫ�`�K���t~q�$�wqm��j?�1��9�C�E��F�)���0�R%�\�> �-v�*'K.w��k^6ք���ڪ��ث��I/���Ȝ۟�:P^�z�$͒ ������Ϟ�a?�oް���	.\���t���l��HMّ���0S~��{�𔤵٤ڕ��Qrsh���'����l#���`!�������<-2h�KD6�YK~4b��vm�t:nh�֒�|�pv�1��^�H����R`4w��\�i<[�C*/m���%�R��mP_X�T�t֣2B��0���`����5>5��A<.��e�t@�Y�J;0�{]N|���ʎC�;����WТ����H�a��Hם�6̒�j�@�;_�OD2�"|/;�a�Hfx�w��|�P� �r�IN�?:K�����]�f)=�v����o�p+C���a���m�Z��vJ�δV�l��V��$�Ƌ�r�����x�P�I�+)��tp�^"8s�.��-�/�������NA�3�xAa]��Uǘ����u�*ʂ�{}������u$�l������D�h��B�pe�����	o.=�O ̀�p;�V#������(�_H����	��WK��m_	zYRAL�~�a���hr�!����H�pIX:h$ga���&��w�5��;����o��@:ia[�}�3|�8^pa�h<|Wށ�0NtH;���|߈ڄ��I��Ѩ����S9��i�W~8�+ȣ�g�V�׳��gO���c.0x�M*(�W%K���jey΅-j# k�p�`gk�~G0t�� ���'�p�b����)	;\�0	�tj��������&��(�����V�tDhp���8��ǜ�)���mM;z��m0���Z8��k?��c���%l��_���ଶ%gP�l��j�<5��� 9L�)�����Rwړ�+��A�R�p����3��G�r�Y ��ۇ�8;�l�m�D[�>��ś��Z�`|�;�����P�L��o: }�?�x�#�{����HsD^�I��j/<��2�w�$*}"�'h�^f�W�!F`-)�2������o�N=��7ıBJ�+A��.(ɱ����c����3��
$��e.��������	ި������� n�y�8s�U1Ct	��y@ ̇��	��vh�-��Z?�\Z)~� =����:��7h��l���7���#yY����<Os���$#�bjn�����1BE�=֨ͳxh%�8���K�Ѭ"}
�OQ5��)�wނSCS�?Dc�-H6�F%5�P`we!���Z��]�cF�J�!M�TЗ�KV�[_<%��G�ɢ�U6q�b�l�N���>�X����eZ�:���,>��D�2�E5�Kr�1��aћ���IY�N�mʶ.1L�����B��&?�5�"j� ��:b�F���W9�-�HN�B��.e�\ߣ%=�-���5�
#�%����.o!j��`a8_�sW��VcAy�^G�w#���
���7�����<��T������;�
)4d�?�W�H�v��b'�Ց6J�j��������hl��I8qJ�r�T`]hy�Ou�OP�LY �Z2�?n�*�z�쌹�'.�������[KwO� ��'�N��Ytw�*Fd�׈�Jƶb4�Y��<�2r/H!��� @��͔o������O=jv	�3�������B~���!��������@JNŉ��n�Xq��E.q�)25u�؉�
~K+�.�R�]� ��mq����\�
"d�v�Bl�B��s9�ͳj�EN����^��
��h��A`LJ�тԊ��Q�����
��Y/�3�v�aٕs������-lK���=9���80����wV-���Y������V�1j��&{�h�������H�~3NtM���R����ʁ�qr�v��U\�HC�۱��_���d��[Z���?9�@yi`8n<IE&�!!*���z�n"9
�goO��N�ӈ��`^����	�i1H�@�*�����̈́(L�ؤ�:���
|�6�#�G8�I�X�Ĝ�.F�ڏ�#� �aG�	�R#������"�P��B�R��)_?KHY|�.���R^��qa���t�����N�H 0[�<�f\o@Ӥ����6-j6��?_H��pS���T��/)[�~"���_lt k�aE��R�2��Z��Y��ĉ3O�x2��n��!�`������!z����dӓ	������WZ@�ǐ��@�e\��/Zʣ|X��s`%̀�X�N;*\?*�gНJt`��hD��3%��;�� ���/�/b�72��*Iehr_SW~\��Z��-�����U�IL���W�;;��;X�KG�X	�)����D��x���T�h�y_*��VkERz�X�жv��HeDx�[A+@9�#�7 M
w�jn/m�n҇�Y�'�B�=���};��f��zx�Hȡ�qF�G%H�Z��j'fN3n�2k�E�<�noK�o�H�0�Wܓ91賨}T*#*s�Y]?s��TL�v�� ݉���(d��6�-r3��9�G�H��~�lqc 0�d�
��Y��k�G��5;������&�g�׽���٘C}�XtL_v%l�����{"q�U�����dڟ)����ѿ�.9��ۇ�)f~��[�O(6��h�ַ�4I�uȽt�#D?�pv��FV:ht��Ły��ͨo�J�O�ĸ�������D~IS���O� �=ǹ�ʽ���ma;� ���p ��p́d8w�L���Zwz�"
�* ���"�h �!b��;�c�Y���^���� I&j��#�wC)kf��2�}w��s���^ �=����F�� �Ui���1�N�(ɉ�*eb2'�d��Rdh�����Bc��o�erk��aYG?.Wo��9��#\N��i�����.2���A�}�k�Y	��9���a�ۃrOJ��5�f*kӫ��Ԍ�HL�u$��ڙad+mr�'ݚ��CR��mr@j8K���|�+�R��L�JH�2*0+�0,~Rg�����iU�4�bUڃ���kr/�n�X���ĩ��V��u5v��@���5���[}j&6���xÙ��iT��P��Z��������'��aߟ0Z�r���v��)�r�4x��N8X����E���a��{��`�c�=������kCa`���}�������2�3�vr��!�Wh�틣�r�{�a��$�<����1V�ֻf������Fg��;�K
R��N�ف>�Y�,����O�Y�~�<B��ɴ��7r-p��`&��j��j8�����V��,_mu� �8\�v|�?:��Ϯ��-dB�� G�P����G>�D�a[J�+�Ml%6c�������	K�ǻ�v�����I/ʲ:�� [{��v��`� ��R�B��!+�T�t�֝�۔C�A� ��>Ļ^��p����v=
ʹ��W�p��>�x�#�{H�J0�Y�!w���_�'��Z�%��z
�����Hd,��p�y^� %�YQ��J|h��Db!���j�i �~����~�.ێ9蛁j[��	$ip�o!T�����/$QS|�j'�t�����9����ƭ_ucT�
D#�_7�Q!�mbsu]H� R��]��U��G�S�a�e�l��.��$A�Y��,y4w��!6��-o6J���!��܍7�.-+;���6���f�ݰ ��S0�sХ|�\�mny�ˠ�I�:Z|;C�2U��+dFCw�!;W���V���9K9ԇ�$�7�1)ߤ|	���v����xN*U�}4`���C��mӠd�O=�H��5�>8�~��ː�;�bð�f��Q��3���u,�^_s[B*��
� ��H
�#)w)h«�'�E�X�΢N�w�x�io����fڻ�H�6�} �[��Iy���=nʌ�yU�IJ�&39i��GD'��k��[4X.Fr<�'�4��T��_|���wV'l8�J�K�kV*�����QXI�b���)�ٲ��$�6*˅�KR�9k�Ɂ���5ܗ��?�6�x˅�[R����/�l[(a^ⱷ�g~y�ֽ&�0tc�@�a��%K9ZLwne'�|�R�mڱ�����5�x{%n'�k�?���ʄ/���p�1,��U��ĨG��Q6q��:N�$gv;6	�Vq�'A�ך��(+7���qyJ��O�D��&�.��+�+8Ɔ�S��̲̑bˬ����p��Q���� 6j�h��3B>'!mx�Lȸ�.���
�e��>�e��
Ǝ��蘆�ӴMz�H��"�R��W�'�
$ #"Dё�,ʆ~�����J����a���JN��P��U�n|%�����m�f�g���(�XݸvBp�GF�uB�ٮjO1��$��\:��_���.yE͈�XV4Rg�֙K�,��T���_�њ���&*
��+ĿH�N�O��V�����xt�G���Y�6�Ik�
{���"�DYϭ2���� '%įT���&�~�g Y�Dk�1��rw� �x��9���fNiD�S^���9x�T^�dR�Ol���&p�����bE 9,h�ϙ�(�ސV!�}��W �B$��Iv�~H�����H*y�uؙK�蘿J߯�u��N;g"���[��@�����-[�����/�r��D�B��{E��e �t�Z���(�u(��-�4��{B���� VRա��P����э�v��#,LP��E� 6c���Õ�#�!5�,�k(��rSϭn���h4��n����E{g�^nb��Z������\	�\5�NM�:?���7��a.D���%�aď�he;������D��r�CW9�A��[��64o�vC��X)�[�>�/n���N<�KޒY���"�-�[�`�`�)�co�5�Z��i_��{*�.�j�8(`�7��6iE�JPN�)��ww��4�
����⡕�K�=��|�8̞�_5��
��h�E �"�"��sޯ >0�l�61B��^^���gҧU�P47�A����#8}>Pbz��ƕ����ͫ�W!�7s�\�?Z�B�ۙ�n�&o8����뵦�N*v�4q�6�	];���T�*�<��[V�r�ق�T��J�A�G\������!����X3�7� �Y�}��4|23P�`N��	��/�Zj��A��j����Ө\%ǅ\NMO��}Q�&n�lq��}p�DB�"�ذ��6G����*��h;�J=3�9�]d~^C��g�K�m����AJ�GqB�C�; ���E��.r�W�pl�Nݞ���Ʌԃ?!�u�a�ٱBn	X�`/pɢ�&��#L���Mptӯ�����6�썞�r���ަl>�O=9݊���Ī�S e*K� �96(|��A�?���,��0��lf��l*��Q��FuYn�eL�s})�Y�@<���B	�jf{iB,�x���Q�s�H^F+d��5����R�0-�KBY�vE0}�E����n��1���N˦�권�e�A]��K['g���EY9�0��bLzK,!	� �?{�%yk��/����l��HZ��"��1['k���7L��ߞz�`ؼ��)C��E���)�1��yv�ӧ'ف,o�]x-���������)�ɟV��X�
��I ��?��ی	�Wx��M`Ԅ#l��2y.��2mgT�.�%&�˷�m��#�Pd��X[�)�d7@c�S���?&W���CJ@8����Ҙ�5�@�BA#��I��|�C<L9�cF/2�̵1���_�Pb&y�E�}��n�3h���g8Ѥf"�� n�;.�}֢�ZZF�����Z$M?5t_ x�tqO�CV��A%�P�h��Ԍ��!�>���zR����Q'��M����!`�Rl�� ��E���?S�C'�#��92ɷ&3�4�����03G��������E";L�G~5�۞c)�M�����6!�Q�y��PG����F.���r,]�޺�i棥�S$������-�9�1R!�P)Mq�p�-$ޡ4c�\�4����N�?��Z����7��MNJ��U�����N=�0$4];�<<����nFz��)���H+��hT��¨\�v�"[�Ȁ���^Z)?j�,�c�����L��U�	��v�JLq#l�����J[C��-ף(sBy�_Q|~��*�t$�7�(VNi�beD�8�B_���D@��˪�S��Z��(m��5ʉ����O!2��t�ib¬�o�Do����0�Z�|RώU�Q`���^�x�a������T�0��3JL8хZ��H����)O��Q�'����P`�Uy�O��8٦��=!�����dֽ!�,�)͐Ԕ؁P�LW����RJ7&�X!8������<�P3�V"S�$S��F������E^K�@�옹K1���H"�	��
zE̔����5���:��[�x=b����!�ޚ���X.P����>LS_tH1��$݌\m�����^?dOK���[�<1\G�$�;��-�U�n�d���]�WDŁ��_[��\���7���ypX��u���y�RF�%?����f���rG�$$���R�U���tHL 1��F��~Ւ�V64�f��v�S���ܥV<��B"0>�ò���5����� M�*��,P%���XK��I��ݟa4A��|!��ޤ7�آ�nD	V�-u�0S1�2V| n��
൱&x��;,CAVJ�uס��Y�ǔ�Tr�w�UǐB9�wtO��ߊ��R&��������>�����_,WY���qmTo��h������@�xtK�Xi(��,�TLYO$��Q&�	;�IfFJ�c�{�z��U*�y^�͠:ci�d��*�Ψ�{�E�����_����o-g��7.N~���A86>�h,���K��c)n�o ���;��%�#��[�5 ����c��a���##��^�ok���R2�6�%��,�"���Pmuu�O�q�m�g�6�F�Nb�������p?��;=���� 
V+1/��3�u��8�ٝyjoӾ�oJ.h�����Ĉ�b�+�pk؈w��J#�\5�.�g�0q#��}ɕ:.���`�bz7�Ӄ��r)+��{=��0�=��@=�r�~�%�Yo����=�Z;�YA^����n9�X$����η1}}�����I���>�	!���_��Z�_
��Đ��fn�Q�kū4pti���^~�k�r��k4��-������[y�WIh6F�����ý���3n����FA���\!/�*�X�gviRF�vymS��#C��ف�a�/��lx�֞z�����%x]�!a�q��F�6��~����]���vX߄d�B�.������wX(� �L)���GLUʅ�pch`v����6	�n�Yݽ�')Z�Y���Jf_8�����X��o~�^B/j��2��}G��<75��M�J���Rp�P�Ts�~����968���?u\�ca�u�7��J������g���C˽�z�����#!��}��HC�m��{�d�Yb���c�	9�A:K���N#�^}���gv[��]�Y��;������N� |D+07�L�c����X�V|��}H������Y��� YӖ=��b�F�8ܣ��8���llN��ptvQ��W�3[�2��|g�q�KʮXn��wF �jI(W�M7^b%��t,eI��Fy�f-��}2���̽�EUƄ�����Lxp-��?�6�I����I�Ԛ^4e�֝mZ��}�m�$i��L?����4��`NܔnY����9;�Ck�{�$Ϯ���3T�XtkL	�W)��E��>�%M1!�Z���W�
s2�bB�Bx�H���^����)��H��uRƹP>���b(�?�l ��D�!�9�_���P[�t!������2�>6�9�7�]�=f�K�[/ϗ�@��
x\��[8�	�B@��ݾ9RH@WRt��b����v��1�~46����d��a��u�� �xˊ�/��++�5�qe��v=E@#�����y33c��H�CS�N2�
�#^���6]�Ō�������t[!��L�Z��YG��;�C���{#�0"d����-�I��1�u���	��*��܁�G�O%$v���\4Od�2�����82˕�d&s�t��@���fT޳b�,A��o�C�u�1��!����[p�`�k֭��9h�I�����`q�4���E=H-z���+*3��&C��u��9����<	r�/��Hp���/_y�,����y^���c<�L_&��o#� d���I#�@�̱�1�&� ��r:C(o�¡vJ[����:��wZ��j (�M� Njh�}�H�i�n����˛	)v�����b��'T�$6F�(�'7���p}xQ���j��n'�;�������խ�Y��r� X��o�]TUKݖ�t�d��롖SR�J�2v�0XV�2�I(r��!��0�1���'��^�Ab��K���\�����((Bl�E��1]��q�1-5�ð}f�7|B︣�}�U�3g@q�P�%���};7w�v[c	��:�)�ɿ��ZL�0V1*��L�x�Op�A��ܫkЭ�*@�Ng���$Q��`g��q�� �n|$�矵�d����s8cJu����{۸�+Y���Gu��_��\��뢅
�0����S�(�g�BS�QX뿉XL/�ۂ ���QY���e���/�dO\򔸖�~oB��TU=5���f�Z:y���X[�-��2%����_������J�?��QL���^ j��\E?��茰9��3B��d7���-�ĳ,eW	$�7����C�ь\:E_���NS9U��}����GIag���7�NT�����TR��c����m%��Vr����jm]����ni��)n�����N�����=ꖢ"o�@�ު�z����z����N
j&�����^>b�Ia�&��$�������w���E�+�qla"#�&ͷ��˫����K3�E:�Ź��^W���_V�z�0(5NxC���=�N��~ӳp�;C#g���|�ENqK�� �̻��t��X�A�o0���v�I��3½sp�7`�Ȋ6�����.AD)�����҅�{���+�H)�1���A�[�#�|�yz��[�O�JQ�9|�L��Ր��/�H��2�/��F'C�[�0��eŶp��@�o%w�+w����U3�aL�hS�Uu�k����:,�B%���<�Si�%�?�G�阚��E��SJ�V?_̍�S�
�)�I������f]gEx��X��t�y}uhY/`�o�ӑ{c����#6�L��iX�����)z�����FB������n�h��+�/j�t�)�A��,��e��53����On����`�
>��4�]=i��K��-~�$ql�[�áQ���f%xv6y"�F?%讔�ŉ#o�EiWk��������	LI�
y�O�Z/������� J�Z��\�*�;Ѯ�`�n��(R�C�)kYc,����6�m� I��7u�sN� Q�����|u3�(m7	9_v�	���3��G�����1� ��8DU`��k��z��G�����r3��-N���HlU�<�	iC= ns�߃Xg<K�9�-? ���8��w�(pI>[a��AY�P\�[΍>'���Ry%�#�>��&O"�;��	�j����Ū��^�y�y~�.@
�X,�DJ��h��Zi�m�KB	$T�I����A�L0�Z	vg%{�f>�=�U�r�vPd�^Gʖ�'1�l[�8��7$e����#��>k]F�,�a��BT;P�OD��9��@���|�ߡ�(fE!�-�S}(�����/� �����:J�˶�ۊ��p�D-���$�1u��>o�a�����	t1WS�H�����ۧ�B�'6aq��D"�x_J���/[���
�Z�G�w�q���q�� ��q�C���Ν�&��!�_���7V��e�����HO����d%�!��&]@�7�n2u�� �:PHi�1,-8�؉*���n���5	�N��þ������D���Ms@¢b��$�����2�{��A�x>%#��"�m�`
{[r��Z����4e��8H���ZVr2q�A:��߭nm��aBj��U1w���)U,'Bv�	�'�֟�z9�Wi����\ �fr��dmU�CS���j./f��чf}�y����YXs�k���I��a�v ��<C�����m!u�N}�՝}�7�3O�
��C�1|�Bk�V8u�,��r��n:��`������Z'�v���~�{ak��k�AA�~z�4�r���4�<E��,h�\��v�%�1���
Ԑ1��k�W{Gr�%�h���$�o����{.�'�fw�$���}0�����9:�@��z�Mgޣ�� f�	[���ܢ8
,c��>��g�	%$L� ���`E��;�nۜ�>�d� ��M��A ��v�k~�g��>	V8���\������d�"��4�gɶ�șR���<����Cgh�;d��qC�*�'�ֺ�� (�;�:�Fׅv�8>I�=��i���~Y�4�@x��J��$D��}�x-i
H�PgY���b>�CV�4sii�F�d�&�۠������D��}�Ap�X�d�>�L6�(���.dyTA6
晸�#,\�yt����O��7s��v_�?``rd��(�'�nzN�STu� %����w�F���Qt|�^T�⌨l�j�:9�m�+Lr}�k���H�bb���<+>`IC�F�X����n4|  ��N�3���I	����_Ϣ���)1��z��3��]������;ј�I�?Qp
����`����(�z~�T�<Q�(5k�e�2�S�Pc�����ia�v�j��)F~LiV���T��}��V�i�-IW���������6���y�G���̀R�
�"�#d�~����Fh�H�
c��e�wZ�6ᚨ[�攛����"�
��_�s���]����+rK�ӹ���d��:�Xh�����A
k�r�`�̀�aQ�Œ�h}f�
��Ě'�+���ԱL2��Fe6�t8m��n�Jr�з90�$;Ï�~7 �k��`α��֛��.aH	,��6e���F�������X�7�$+��9��ץ��r04���g��4�|I�_�M��j�� Ħ` ����b���H#3���<���+�7����С+��X�c`�85>�Ss7Mf&cs�`��;����*��T�m�R���5Ü:}ʗ�6���ٟ���	���j�f���W6E_9i�/��FS��]�	U�IMiNd%o�;ZA���Q�P��I��x2����1����:Ap�P9��sg��Aלٙ�]���������4��9�8��E4�$��d��@�ج�Tݷ�ţq�#e��BQ��C�ź�#(]��FX輵�.�7B��5�~��߸J��$XJ*5]�ι+�?^��ő��-"C�q�n�e���B/��\�sc��0Τ�LOS��ݛu�����
��%lt&��^\�X�5ӷ��t,�������Ua�j�7�n�b>R�I���&H�Ҹ��dDX@w!%�8�X���B�R��{�y���U��f�TɈ�g8f�M*�%�=h����%C��JB�B��G���muI;������*+k6$�Y�1��@�HDNԕ��/L�\f��^��xSLv �>�&���<��!s�1�Lb4��� h�(�2�C�7,���:�Z�O�$��:�ũ��Xk�o���#���v��.+)?~C`"������X���|y��IGۤei���5x< 2�g��x�i�3�J6�pή��65�&8��h���H�
���-5�aQ�k�eW@r�B���%�{H��dߎ�N��T���:��5��ԏ�7γ`א�VS@`X��������<W�*0�eC����r������/�<�
(G|(���vUp;l�W�E�U�+5|dVͩ�.�b8��:�A0��NB�,��)��Pe0Fc�/3���~+y��EN��)7�;YSڶvL�f�B���T ��e�G�D�'�=2��?�{�ޘ���_
`�Qg��|��h]�$�������t�2*� �O��yOm�uLG�M���VlIRP��Gfr����"h��a�_cNY�]��G�>��M��LP�ߔ@�op��՚h%}��BAď5�{�d���aV�۾��W�ON��=֡��)[�ӷ���WNO0���w�w���Q@��p���a����@������ʘ���p4���<z@
I��D@�Hڱ��Gx��4���U0���o�9��yjxK���</	�+�Ba�":dB5b�y=�1ȧk��Y���Y_$M���xH���b�3�BR�J0u}���� ن��`�h%iĀ���ּ�%��C�鄗&�pD4-%Y�)��׻@��夦��#2����؝ "x=]�"2{G������Y�G|e�A�(sŢ��^|����ˆ8	��D�V6�|^E��W5jaF��!S8w�YH��t8��@x~|�֫�'"�,BE����� ��kiej(St(��$����eֆ�jS����γ\���M�� ̪i��t�]K@y3z`�o�38Q� �?����Ĵ��\�  n!��z�b����aE7$k�ݧ���Wv��{}�F���gZ�?q��44��?�B��^��� C鮫�s��ҡ��6�t|�����C�l���f�e4|���m�A���?.���DM�IU�Ghg��ݞ�q1����`���+<t��+CkM6��=1��V/ܗu�^|}'�m��C��v,7$�<B�/�r��K�].g�A�2�g5�>ʩ��H��w��������7���`�"�|�⭅6�Ǭ{�5흌���O@�
-?�Vq�Wť��I�w/�����Xl:��02�8񩂐�B$��x� ᡡ��1�ߝ��E{��p�g������+�,*X�k9k�v?t֘���m��e��3+���f�oeNDs(�O7{��j�����P1m�|��r�+g~��>��+\�&ȟ��
"��->�҃��>�[E��'�'�x]�5r1��FjI��8#VI��І�7���_�
�"8�,w3w$�����K�U)�h��H?<�Ԩ2nN�a�;D� Ϙ_��&�nǙ����v<�ٰ$��4`�U��B۟�ʧ#I�8��me��d�eɃ��aHq����� 8i���K�P���~B���ĸ+�r;���=Nھ�:�ڂ��b��� �!~��c�7`���b>z=W��x�3^t�<��f�����柛Ў|̤����{��%U�sP����D��a��PN����<�(v��A�`߅Ӹ� �e�x�wm>4U��S�j��Dծ8�� 9�U��d�x@e�"#Q���*���t�3��D�BC�և���B"������K��=&�'�Q�*�4Fw�E8�(���C0*���[I6���Y��xi�[yD.�*K�f�s����uXN�{g̨��J\/��I+^��QI��7���n`�blk`���R��>W̬w>y1@����s�-I�1'D��-/����R��&��6�@�-dj���Tr,���\����A�ɻБ�݋�?#d�������A"t�j�oLLM1�4/���D��$�����{q�N�֦�:�6��E֬������\�ؖ��l����AIK Tf�]8��w���M�$Ќ}b�<��sH9�=����e�@&��q�K���ȍ�GC�D����L����\�l1X�O���t��֍��)�#�M~��_�@��K+��o2��ߋ�U7Y�Gv�(ڒ��O�_F�O��q�����D?ٰ4C�ud�Ga�I6�V�t�˺�M��pt�	���(������&�^�ܛf�^�}!�N���k�`�t��mK���?.����i�2��5iju��i�;��i5�юM �/�W�m�P�N��)��U*b��)�%�:��yی�a�[�UEm�ɀ�E/5�BG�/
8���ݨ�I�;�c%o��I��x�kM��~�jkR���R�U�V�n3�!��܎[5�Jz�F�o��$%�o[�;j|��*�0�;.�h�ٓȎ)>���
݌C����羃a�z���%�g��rG��c|l*��Ϙ�&�%Oą;�6�_f��1��u�\w4���5˭��N4��}����d�	3?W%�{_���!�~���#����{�p}��2�K�;��`Ȝx(���9�k��:��3�<���;��y� Ÿ� ai�7ݴ�|v �>��y;�Y�VZ��j*�aQ]Y ~���QV^�2�[�lvQ�βu�d��[^>���\M�Fv��i��&q	�6�~�����4SKp�>^Bt1�6	��IH�4��tp:]��/�M��WH9g�L�$9�E��d���~ʌ�M�A��er�����f�l��ѻ�;%(p���ބPv;���z�d�.f�;���L)E�6~����s�M�r�2��q%0��K�&�����1P �Çz������2�aH��LU��)�Y��a)
T�������������U@]Ώ��of��uB������O�y��U��v|`t������85jQ�v'~ʠ$�[�3'�r�Y˱�.yr��x���0WĽyJ�
�`N_��(�����ⱦ��R$��D�;A������!4Q�)(�����w�T��3�c(�L�[�G�t�W�"*�^����Y��dH�K�{%&��j{��E�Z�,��W�3�"�d`�_�,+#�����Ls�K��7<���@!l�80�Qǯ�<?��T`�7¶/����Q(��j�ީ��\t�,+z��)��Rc����~/���q���E�"
��=��8�8����Я�~��w���Z���(�\ ����o�
�[���ϧ2��6���#���I*\��M`1әܲ��=V�Bg����6Z��A'�8��V�s:�1�x�N.Ǵi��ֲ/�h���,}'���;���N-��H2�%��	��=)���kv>��b�^�*�E�!�O6�;n9�z� �>~^�T xJ9m� ���E�����v��w�vpB&jy)݋��mܵ�"�t�A3h��|0=ޢꌕ��x%�V����AE]�6f|t�h�q6\k�����x�W�:ƚ>������ 6�#����|bW�����,5/�#�H���}���*���oؤ�!G!-��cZ�J,4�q��~�)�5�s�\T��0#�	H���s�x)������(z,�ؒ#�M���e:~c&ݶ���*����y�J����h=ap���
�Y�M۬���?���*#H���^�,]A\�g�\����NH�e.+�גxS�bX�;��-�ҫ.�qC�!'2�[H
Cw�q�2�`d���%��F���-�5�qh��Vv��gv� �7�j�n#yeڶA��$E�����Փ/�]<�>��K�� ;X��xU��m�Җ�>�5�"��ao����3��X��Y��V��[�5H8�<��)�c����Ѣ�SG��z�0����A�U���v�]�;�O
��&�!��Wk f�JRXS��&�8u��S�~3l�a�7h( T�?��3.�b�C�2I�rH�ݐ;`�,�Π/m��O���&H떺�F)6I�]Xhw1�v�+��f��&��f�ӟ�tcũ[�z�l���7ks&z*:�El��� �o�����&�XD�4��;�� +{����3@
ڕr��á�1�U׆?���T�*Z����7$�!o��h�#�������,�� 
gƼ�jg�?�x֑�_��]t��oG��]�v�$�qlB�@��?��T�f9�^Q]����`J�}��"�J�tϿ���Qf�2ΔPIY5��+�ߎd<�lY8B����oe�)ѫkB�d��`��I���W�YSfiX/WA�SmB*� dV�&�b��q/�����h���)�� ���
:�,���L��,ٕ��S�׹�eAF��zTt�DN��1�����h�K��s�l��UJz��>��v����*�H�%k֘���=���۝exm��NNu���r;�R����q������hL �����\�&��8D���M��dLmvȻzqL⼝���Q�}	��h�c?��3�g�X�y�p0��Ejԝ��5��lVT'N�g�N,��C���e6������^����j-w�)�&d�7MT�� u���/N��H\D��]�vHd��4�7��=J.�]���L�t�ƚ�IZ ��	qt��X�kg��^[��x��.p��v
ԛ��� sqN*p���f�&��T �����ˑ�ml�4.�6?��g��[�
�)��;�ұ����f��	ѯv��nf�������;�P*8���919e�S-y�);y!�[@*JyM�.�sml���Hi�[�Εh�PӋ�̡n륅���ASNv>�cm����ͬ�5S��u��nER�! (���R�T�Z��^^I.ME�bzj���R�E���*��k��:\�R?�6�B����@sNa��``���{.�1��c��h�9.T��/Hdq���Lk7� �񍡦�j�X~0F�(qc��.�'��(���(���[�:���G����|�F�Ļ=��m��j��7���0�w'��(��G<��X�k�5Q��������h�K��]��Ӌ�^ŕ(��;����rZ��e�Y<bP���5Cp:�}T��K�L�:�W��7�w&WlM�h��R�m
~�������V��v}=R=����[�+W�3����e�W�b1����J����v[�>jO�X�ve}���8�c���{�&��X_��\��y�{�X+�Cy=�$�#�΅~mg	0��IWQ�ax������
�P�N%�"��!D�
; ��l}@�2�ׂ�66��&F\b����(]��{0)U=��s�-d&�G�R�8�4�A�&�Y!'�"vxZ����R���,���cU��h�;�g �FtzN��蒽Y� �ȪtV�{~�@D.'�)E,ܭ�L0�GW9!W��t*�2iN�~J��$U���e<ͪ�?��*;n�c��k
f�-��w�S9�L@x4��+��n���)��I�G��KV�(g��n�d�c��<���m��4��2��>"��y48�^�|��V;Т6,Q]e���Z�MP�#NЧ	��0N�ԁ_3A����m�,�p��2&;�m��Z�v�L�C���+�;�-��gY�'ep}�>zoɓ=�M�7���ߢ@�ڙd&y�s�A����Y����(���v����<B�(n��#*M�rB�o,���f|>I#4�^���d��kvj<���Fiy��(2�a`�to��Ex�9>��N�Zr��^\rs����B���="�
({8���i�j����~��T���3�n�"ю��6A��W3�s�����*�P9"J<?+�1b�ϥ�K��_Qi槼=Ò���7U�r.���Ӎb��XǴoa�js�ɗ"O&7�#QrA�/B��R���1F;볾p�Y�N�#�����"�@�2��H\�� n��o����nF�����[�\]���@O�����#@�JOI��i����h&xt6x�ɔ8��*���8��+~���/�����oʁ�F0Zh�YK�J��:��J��@���7aԣ��)�P���C���yF��/w���3�F.[�\��tf�Y�%$g�݋��U�X�'8S�w<�+�%%5
�g��I��qo=>D2�>�O��J+��M/��4H��k͑^1�?� �d��dN�{�J�y1t5�̀P������z�&3t��*v�a�V�
�)�F7uo7,�:]��5rѓ�V�c/FЧ������'�뜫L�<�h�4���ɦ�����B�r����v?������sU�J�ĕ�t��N� 1����� Y-��5#h��b�$9��}��b��Ty@�X��aL^�6�VC�|�����p��UAs��r��N%�{o'�I������X�ugH�U�_�˓\��/����g;Ŋ�C#@�*�����CBc~.��Me��2ce�<���ؼίKH�F"���H���B��b�,z��j���%'��Ⱥ������dǐg_�}�v�F=����Hr�]B�{�~�{�jY2{±����9���UE���"1i�tl���,���-+�,;�f',�5z<�M���$m!+�u=}T̃����o�G��7,�Z�A�(v�q"���z.�~$�
�Y��j��.Q����Xl|Udcy5�/&�#.D��FxX��df�3F@'�/�U7�z<
�I�J�`�z]���{!���&��v����=qtu�v�Gf{�&��L���d\���>������S;/�/ؒ�Q�0C��߳�:�Α1�"�D�i:��.�ɞ�@k�1Eׅ-��9����'=}��g�W��o�>D`�ȥT#�����3\K���ժ��Sw�\}.HV��l�{ߘ����������e�Ӭ��-僭��ͽ=��,G�:�^e�l$Br�~\X0~�F��C�jY
$]���+<X�np7cnV��N����m��I�;X�~}�&"^�(��?-�{�����@�Z*��{5dk��	�[ڴ�@���y�r�(�0�k��8$K�Q�^w/�B�l(>��*˯*b���x�/���^	�7c����q;0�,;�5��c򷆠ce=����,hi�-Yd�u��m_��b�2��s�-$d� R����[��JZ�.R�S%)�R��ϸ�� n*��u ��{�Ͽ�m8<?�h�Z��9�q�h�[��aD�蚝����u�ޣ'r�-�4��=��ω*����v��ߕ$g��S"�$@�D��Ԏ�B��Z`�2�����/��S{T |��B^���o��8�p��/3�"z�E�IM�!E,������=��k;�I���a�J��5�s�ny$`l^���2
-���Sݐ�OH�t��\����
�Y-�H���R�c��X��%F�0�s0Q��KduL�*Q��u�/�#���SUQbY��wc�Yڸ(p�!!Ն�o�mP4�ە_��Xף��i�H'_k�$���?�&�	-�,0���(޹z��!Vy�^ XWl���������˿�� ��hokOH�d�׾�g���Ṵ�*�����jx��ϙ�ɶ�/�%X��a%�XG6 �c�;�Y��(�dkƃ��I��Ћ���a���i�}�L�����Dv7�!l�=�cY�k��x1����cM�
?�5�Wa7�wDJ���jXs^�e}E���6��hD�x )�?OZ�@�m#q8�
�a��ounh���E�b��6\ܮJ����L��f��)N8�-�4���������K�O��������u���sc2u̢�뉚xd9�⤀��$.u����UM$�����U&��/�#�'K�%�X ��)��ohb�g��5���Ѓ�����8��D�c����mh{��8��ȘyVz@g��7��D�M�K�S�R.�Q��I��Ƹ�age� N��{IĸG�"7�/� i�4)�dJF�"<>�Zꉶ��1����~���O%P'[��_��Gj�ܩ�z�H	�ę�v��Jfa�a�Q��e�/�#Zܹz����X"��0��憄�YFp8��-2�t
M񲬇ꋄ?��(�q0œ��L֠�Ţw4�n��&J��3�_��n��uo�Ѝ����I�	Y�}*�5c�l���`�zU����4� �:=`7� ��|@Ǯ���ʾ"p�9,��K9(3��fcug�&��S���RCZY���B;%|Wz][_&���#�����n��*p)��uodߧ�YL��lBtN�$���U�e�᤯b[�a�;�0���j�8��H����sv�� �1$�"�#
0m_�=[�F{��i�����6`������c�{����z��T�
u��+��������u-1����0�S1^��9�A,�vwI�34:=�J�<���Z|����Ǒ�dC<���?�i�X���XY��u��Sibot,K��g�׳�)��H�93˰�F{aR�����	����fޮ�ފ����nQ�rzy���:E#T�D�u��}�uy3|�q7��h臶�Y�7����p�B@b�}�:Q?��ؼF�X@�OM��:k��m�ٟi�M���8�n=Ƭ>�N4�d�& �T}��ܽۿF3>��s��e�kO|�:����%L ��ı�2��]�Щ��i�]�穝x)F���$Ͷ:���H���M�z��ޚ�J@F�J�t���WX�W�����o��*5{?�Z/�n�?�5��okzX(%�ٞ,Ս�4?�p��ŋ�Å��W��mU����鮲���UHW���UJ�����,�qb����)-ή,B�J���'��+�k�`��جѝΛ;!�U�k>#��:��
��	�Ƶ�)��o,��L�]i�20�!*ݾ��F���ic� �G��C�y0�T�y��e/j�� U�V� �W�;ע������m�s���/w��%O�&��U�gэ�a��\��4�>���"�4�Y����`(����U7�T��Gۻ�˅qX}�6M`�(���`TjU�'~f_+w��a��!�*^d�$���[PӢ#�L��������]/MJM�i�Lřq�`eϱ/����;iq�D��u=a���x8"�L]��%�Tr6��Oq2���y�~B�x���Y�U�F�Ε-�
��C�-��W۽-Y�i��т��FN���(?=34a�kQ�����*�v�2�	{h~�� ��H|x~6d����Zf��i@0n���<��r��$^��Z*!{U�F٣Y'�ֵ3�9v���d���z/t�����X5��*W�{�/'�2&p]Rq�,-dO�Ldz�C��9���B0�N�(�u��s(W��b��ɉ���0?_�_�O�(�1͹�㍉���-oL� ���z�^���c���y0y�Yl,*/�̃?�t�xԡ݇H�q���l�WF�vt��vhK�W���aI�2q�Ʃz�A�������]>7d8�nr�B�ÒeCiIm�vFx���p$�����S�='���}|-|�Z����x��1�w�:rG7����]�p�Z��t�I,ٷ��"zm�#2�,��=�	&�@���j�#}7��s/��b�C�b6�l�ߝįiJ�ދ���^��� =߫Sh���� <�^m�&�l�g��wIu������<�~ڧ�6���`�U��/��}����pXri�����	tt
�i�;��ޒ�q�."A�
D�l2�����B�<���Tsp=��h�h{3\�fve�U���a����)��Sv���&>����|P1n�d��PBc��*� '�m.���w��֝J4�8>E'-UB-�c���h���ǭB��v}a�s�G�hc%{E4!�,�������-���]�LzB0��ڐM_�A�U����6�W8|S�s��r�^O
���7�ꍁ��%���ٚ|�C�ǅ�h#�\�N�v���e�s(ټ/)b�v8H�$�ת_x.�4� lڄ �'�8���Z��&v\��7[]��:�,�A�
:��R�0��۔Ͼ�wI+�C�X��u�>�K$Ư��xһn�N��M�r��c�Z�ZS�Q���^�^�ҹ��e�(h`�W})�_颔�py:c\�K�gMW=ը��Gt��;ɓ;y9�^+6͂,O��� 2��S,A�$���XC�cs���l:�^�f��{��h!��t�����Bt�c֤�*rH}�K�v��kl�Os4�����퇠��l�x9Qf��ӇؕE-�Z��6d��� >�п{Ø�t7b3�M DE���$s1-]f���q�
%~��IY0����@�^iq:c�;�U��8��qL˿6��?+pY�ש�]3G��̞��,U"��Z=!�_ H~�QL�)�� ��$I�[��Vuʊ�he��z�f�#���������h��#/�1"'#?4��6�p�UP��Xٛ�b�Ib�z���ۀ��8����LX���[���)eFW}	*'�6�{����$S��@�pR�6j������>��3a�l��J�^3�L1�����l~�]c�7�`,��HM�u�mcp���3�4'm6��ts��ҥ�?�'�x�6K*�7��;՗C,��$�����<�[\�~Te���8��L�G���/�S��w�Hk�����h��%��tr*}kb4/Wu8V�`�J�����zhE�k}���6!��t������;�����윗ͺl�I��N#��B��F����C3�>�n�I�;.����d�f�#���)�0.���Wk1;���s�H~�9Ge������m��Wc����x��Z����軱rS]�����{�h�ꈎ:N�;�-�T�'S�@wħ�i�=B�k���	�tr>Bfwv)�6��7GA���MYoB
��wL���m܆,�XK�؁S�OC�e�)�C���:���6Z>48�9c�X�R\��#��%��KW]�\/��Yy��+��&�_5p�Y���l��	�g�,,�=DsC�:+ �w��=�����e�Q|�2�f<���s#q�,s~����e"k4+�͊�von�"P]��D��5���?���=��m�hɞ4��:4�/�5�"��6yX�V�`b��m�
E�#1��9��!�S��E,ݏ"�sR�>�-��9�B_ÿH��C訹P����<���>�Jz�vߡ�	��ȌP0�.Ʉ�[�{�L�ou�%	�?��A�{�s��ч!P����J�o���^� =��|�+V�4%��s2g� �� &�X���D-K.�jC�ї�hä�h	%�y��<�Fc,m�
*����k�?�M��@���KI�F [�XR�͌���~��Z��R�%�H��e���?&}ܡ�������P7��`U����������;(h��S<� "��|�i<�x�ѝO�\�%�H�De��_I��~""e��1Z�8��\�(j���T���}"_��+�W��f;�z��3WK�(�\UG�M�����
�-�$(_ʻ��S�/�����T��q��
�%է]�����d(�r��{��1�c���l"��}�ԮukG��+赴�;@pÇ��9�DW$޺���YpAZ�1�3��/�*�\;(��3���4�d�:��L숦^I������:>E��j��9����vʗ,!ބZϰ�/����=��z��j#Q��6��J�8&��
��N��B�zT�ܳ
�,Í��\�ۛ5�Z(��*aT�ᨭ�k�,���.��N�,�;���"�`�T�_	���ݼw��i�d�}_��\菚�aH��a�:����@u(3	�V݂e�U���{\.�� Kkx�l	g/n�pk�4o�$�G-�!0�1�ģŕm"��F��'��]�;������[?��Y�,�/RIw��G�j����goS�Q�a��ﭔ?,z�q��lZ���̨��UB�YZZ�ͼDe�Q�1y��,�여!�"�VL�&��q�-F`�?s ��ύ�)
�yq�8HlD�v��w��n�����J@cȵ����[*z�R���n
ׅ�4��YX�'�b�%Nnb��%��d��V�n�@"4�u��z���;g���S�0m\��I����Ien���xp��8��E}�@�<��	F	�d����vJ�Ū*͗�G���W.׿`����a4�g�*���`R�JB�B�1�ό�&h��S��D�A�O�
@F� ���@\����L��o?�mf�K��q�_A�*+gj�M�D��U͖��X�dTHwɶ��Y��sX�~j��N�H�:���-�Ю���g�����T���D���j��W��0�S���LJ0|q�tP��E���(6��?\@-d�S m-�3vz5�W4^{C&\�{�X�ڑ#������l��v�� "�b�
FWB�skc荬�OW�	"^j����k35}]�:N_\T�`�m�)�C��CUᑯ�h�Z�r'�܀F�R���C��)���e+r����(fu�]<��!�~�Y���j~�(���Kz��[t�N��He6Rq�9� ׀����������%
iN�=���9�ᨑK�f��z̃�]��E��lB�����\M�`�|x���{قg�SE�:����?p��Z_��x��Du����;�z���ir�"����������ʀ
�T���2�P��aX_p��ә�����㒁�#>+�Ռ��˪"r��T�6r'ԍ9�`�bEba���f����sais.j��<wP�����E�M���uz�tQ�q5[���X&M�#�_|�q=�6�|��(#��
�������h-�@��74Ob
�|�v)kT��Z��e~�i�״6qm�V����?6��,� R{�����ՆT!����M˦#���G��p�:|t=��l��>Y����[��?�d�S�W��!уcz��.��.�I�W���7�E̲~�RP*(x����W�����MHîɪu/T|=��]]e�����*#�e*z��Ǌ���W~h��U���M �8m�@;�޻-(����S���}�@+&[7�"c}j������7Vd�]C��-��ﳈ� �|�by�|i�B���u����@���N��=?�B�a߷�T8dX���}f���q	k�&5U��J�WX�d�u"c�uZ ��F�&��eC3O���+��kO�&W��h7����=r��EjJ����9 &����.H h)T�����'i��r�?X��w�4��l��;�D��d�RԬ��\*�'��?
΀�T[sV5�諡ew���8v�M���KF�GxP���a�ER͖��v1�%���g� ��e��H�`V�����N	���Q�b�\f��}��X�j�!R��(�Z�f�O6�����%N�<Q��!��ձ�����ۉD;����=�*o=�U���=�r�^�=�%&�<����j1�$��@�{J�z圲O:���h�UfȌ���.��g|���(��e�6���� �,p��gg;���ao���|�v�J7�};Mvf'���}|�ʴ�%�]�b �I`J�U��ɯ�/�����\�s8O�L?�N���=(�X4T���w��$!8ۘ�9q�`KDH|Βp�(�F���$7 J�ֶ-?Iaz����J�s�D{CL���f��;BS������nG�ZqtF�D�*�}�u][�a؉Җ��d��+�����ݗ�p:�w%a�h5*�C��a����Q�JDY'�Gs�����v~�#FU�k0J!�a�3&��߱��-o�?
�2�s����3(���r��K��X[��ϰD���҅�I��	*����ý?���|vD���X?<�����[��]�+d�o�����/g��;�x��+b��ܣ��ZmV�ǏT���ė�~�MɠEe�������Ŝvڊ�n>�]Z�]�^��k��9���5�������������G�M�$>>޵���+"�>ܧ��y��p�2����ʚ��������h�Z^��K������@�3`o�c��ӒW@=#ǔ��E��eu;Bb��j j
��A��X?P��3s9X�I��z��^�`&عu�Cƨ^��E�;�6�ҧfX-��ػIӿ�U��W)���G����CY^<T��;Ϋ�c���70{)J�oN�&X�x��*;�~���+�b?I����un<�}$Y�Rj9z��}%=߈������eOh"��G�h�{�̪�.Qfh���`���d/�X�uD3�H�I�m
_��>x��6tʞ���B������B�S����>д��j��<%cY�_Y��g�J�������*ˠ>'�gٖ\x�t��s$phѫ���t&|I,���!]tQ�r�d}O�1���co��(Ҳ�L �u��1���ga�C	0	��A�W!���I;��	R	v�%�x���}i�TРr��ƻ'�8�Z8uL�*Vv6el��J t���5�k��?*���X�WmW۾����O�����g��2]"�I���žՁ���6MıxH<�>�S	>�@�-�P*JJD�)$����������������C�$U	�$0��Dyg�聣
U��v�<i*�mK��D5�vp[#JZ����ct���EH��CˡY�'����*@�,l3i���	=�3Z�K�/�"~���6-��%Or;�)G������4��}��d���
6��S�p���Eo;<��^c~����Ț)E�3�-�c%Uf��7��������YF����a�g7�AN��'��GsT&���p�Lض����'[�����a#�8��T�Ǩ��e���֊���g����@A��B�z��t �t�>-z��R<����i4dM�L+ő3���x��An��)˵|Bj)*}�P����kW(.鞧��xEZ��������<|b9��߬g�h��K3;���L(���h�͍V��mu���s���}%��=��^�ế�[6�����)��c$������G�Qm�SLx�z��ӡV��(����u`p�<�B%�spAd�b�;�b�jӟ���a�k��wEɝ ���\����ѰA}�?�ˋcD"���Y�O���3��B� ���Pt�����^��L�I3|9L�/�(mB�2���x����{ƪ�
U�'dh���$�%�����
:��W�n>��HIe ���*���g%20i�G�3�T^B�U�Ҵ��~w�h4
�djK贔z�� *��X�E⠟T/6?St͵�S�ؙ��n��:/�t�
x��en숅��t�N,؅�(����g����.
��V~(_�`��Ϋ!��
<[�w�,8���8�s-K)������S/�A�$�����ä�h�K�Zcym���D�F�8�!/uT��y��@�T+Z�����nǦn�z�0�\cA��K��`g�TrGEL>	j5˩��z:�V*��w,�M���	*��e0*��k�="Vy�غ���y�/(b���@R���ʇ��9�a��K	�}È���`l:��퉾�Yp[�?����aNω��C��S̃}�ŗ����:�P";������W_3�O�+��9q��s-s�f<�O�d�wB+CU��Ğ�;n�<�k��\�$Н���%i�1f)� �+����ϙ�vP*� u0=^�%���H������ J�M_0V�ɶ�@7�E�t?Ny6q$�v���"�R�6<钇P߬ξ��ON(ƕ{8��iY.�<͠X�7x� +1j�s���D��G��u��>i̕��2%�ڄC�z���I}Hp�*`3y��c�S��${��u��M��;�y�h7�XMc!�E~ӞXql�#��V���yA�o���W��O��z�"�l�̻z��-�J��\<t�+}{Ǔ��S=�.Z��0Bΐ1�6O�#�=�1�9�K�đ�*!E��x�%�G��qK�f�P;^����`
i
D� }��}Аdt30KZq��q�"�ƺ_E����H	:�<S5|&TO�#��\�є��AuY�駋D�9υ�9�T��p��N�T��nKv�u��pT�*X��M��و�D>��g�Ԏ�'�����e�W=:��<U��rh�\p�E�|��*���0���f�)��������)����&+{i1���?Eq[���f;�zZ���T\7�_38�8���LD|�6"��ŃKΫ�tF0+|VT�!�I,?9�w�ε�XS�Q�h0=[>�~�{����֪��B�A�ʮ󥜿�RE���3KR4(x�h��?�bb{ɗ�O�F�u��L�'Y�ǐ�T�S(���X��_~G��VO�17<�<��s:>�P�K�>�:��v"��QA{d�������`�UT}@�s)pQ��|P�����ʙ<EPm�������5(�9f��T~�1wl�:��{s�|��D
�db���qj��N�ʯ����E8a��\0NN�om �<}��AU��=��O�����0�;9#\�i�<A�=��ri<�+�e+J� 3>T��R���X;�}�'�ǁ=������$�����+�v2�AZ��R������QMv�E�=�g��`�/�e���Z�ʉ4�i�\�Z��\���^ǁ(�h
��Q	i�_�{Ls����fʅ���������n��_Ǻ`!��,���o
v�0�tpo&�e-��L(+_��cN��C��%#8��{!���l$�<:����l.�a��m�������<O�i����8��<��������H�)B����|V� *33���]����&�� 1��,��nB9�ȵ���%Q;y�(R=V�A���l��}�6g�4z�v.ڴt&�z�����
*~��������"|��mT�v����F5i����)n�&���3Mp�k<�5�TʤD�}�Ϟ}����xΔa�C���?Qp�.�ᒡa�������:�+�,�x�����RN��$Ǭ�[�D��s90b��:��;��[maN�:Y��#�!��Ch�wv�/�!�;')�ST�п�q���ȫU+a%��6`%D�g�4Y�=��G.w���uHLy����w3
u�4�K�X�8�-Ѫէ��ٖ�8k�Rn1��,k�O]���5wYPo�+�V�W���SىN�bj��߳u��0���oLh�D�	�0X,CQ�Fe��ɵ-ϲ`��U�)�un����}ON���P���T@\c�>���Uo��0II+��k��DJ4��xh��a��Q����@� ��Gg���~���V��:Z`�-�4����koA�{�=���R�0G��	ߊYUoqi�����A�{�)�''����LJ������Ҁ��s�Ś�ǆ9��+�${����Ɛ��.<�D�O��� ����y����\�����9ʂPK#t��|z&W]��K*'����(��]]:�K���﬩�(¥�ʄ7�v_E��O2'��v����"�����92�)�m����=�2��ٳ^�B�{WG�З��[��
�^����������i�M�� ��/{�1���+�<�Mv���YG�K'���2S�=S��@Y��2��n��"r����7��T����X�=G�Z���Q��B���8a�#�|ό�{$a-�v0��k��8u�k���6�K�u�2>Ƕ8w��\�+���4D�
ql��Hik;���RDXRK2�Q�m�
��T3\$g?�ߦ{�sF�W^���yg�+��pS��=��4\��S�$�M�ƽ�(�A0*��M$;c���n0�so�*��Eڛ0�#�T��tB�\�t�ps�?��8~�Uk�� ����u��#PZo��H�3����2|�"��-�¡;w��1�*��v��n}D�5��@o�_,�����9*7v�օ!�	�p'Ճ���:ͼX��/�`��SM�Ze,Kmb�~`�1X�B�t P2���	+��PRAo�3;�?�}�y��[Hc7�&4z�mR��K~Sd�/\S	E'�*x�V�8�q������b�t�F���B�V ;�״����~��F�6Cس��k3,2ͫz��x�Q�-VD2L��/[�$<̄�}	�C��CRJ��6!�����AR���3�L�fC�afZ���H�қ�������ƿ����K��x4���j��tm#�||Թ�|$O~}M�i��I��Fj���Tk5�Ɓ~ơ�7��A���a32�-i"�K�''��,�nm�;K�DM�,�U�e�C�f�!G���c@�Q&	��&N������8��#�� p��>�P�e7p,6�?s����Iv� ���ufDZ	���G����'HT������X+�r�D{����. !�}V!T1*��n���R�t���vz�vJLv�[�bw@�#�:��X��g���`C�?�bG<^i����b!i��m�^6Q��T���	�ў���YC��O����y��:��hr�	�N�E��V�oO�+�@o>��)�w8 ��p�,������FU^�yM�+�E�{a��� ժ�"J ��(y�A)L`E�$.w_qp3�Z^�Q��4�D��\�m�2k�i��|<7���" ��񋛲B!�W1��\�,E>�7����$_�	tɷ��α%]��9���$!�G٨� ;�@���,ڨKݒ(mw�F��yV5p����_Z���Pܵ<�*�8 �'Ⱦ<�c*���մ��i#��/�=��8��<%�3�l� �;a�����2~��ʤ�}�P��� pӅ`��3d�õ����dW��9�U:��2HC�!F��`BPϖ�(�f<�(J]�D����Y}�O��!��{Y0��5�N3�8^��M�[GQF�ƃ��O�ѝ>j/}�3y�I�	7b�7r��ņInkq-6��Z�,ZALO-���顦*���$BɎV�Y�������J!WA`��:Ѿ���V_�2c���e4��it� ���1{^;�2m}��X��7� #���u.Ljl0���ƈ{08�)VS ��c[�4�.���rݵ���(AI䈋��b���f4H��w3z�Cz�:oh�&U�[�T���)�>����3A4x|Cح���)��.�(V���T?*{p*.�F�cπ�X�n�k��'W�W2�F�ju\5q�A*}��O"5�U���� ď [�to�6��>��A_Τ�kR�&쭔R�@;dڒ�Wu�_u5��|�m�)��OX�s&Su�@������xk�rűA۟®2�b39�S�d���z2�B�ؽ����}!^B��!&!HE\
��v�tF\�Ʃ�Q Yĩ*�d�j��]ꌓ�qF�Q��q@ϧv��=��ʎ7�a$
��۵��YYC4\�-
��50�*�so�F!��:����Eg_,$�ri>���f<T�읠�Hz�����WyW#e�HT?�$$g���p�|�ZAI���q�+<�2t� �Q�����+Z&�L�ߣ�A~G4�!�Yg�6����=Kt��]����n�X����W%���>_|َ
v��I7)TrM���Z�K��su��ؗ>w<L�c\9�����ν�J��Ꝙ,ɼ�(

3�te�2t�tW�v�I-�CG!��L�U��2�Fը���*\� ��T*��ыQ���=�Q���{r���
�ҨQq�*G���킅��k�Ny^�۫MؒjAqɎ�4'��t�~�K���������ق�+s�V',����GÀ�#{1`ɿ̫W٩��y4/=`��[zp�
ĨS�EB�g;F��ʓp�
�d�*c�2.���g9�A<Ӎ(�iX#�&{[\ =f���6�~O�'I2������oQ؊��t����c�e6����D�e)7=g?�✦;,��+�V<1�����^�~��G��;y.���i��i��Dԋ�h���[V��T��)���3�K<��pot`W��/��#l1K:���./�Eo�%0 ��\��[!�v�Չh��P�H������ǝ�3��)�&Uf[�/�T}�8Ye�C���a���oY+y��`�w>G�փns��k;�f�����a��e�Ȼ�J9 �@T��X�t ���Y)�	frNI���FM`	CEp��(�x�߯��0 0����c+�Nv����Z��iҲ�<Nj(AS�����vZ��N�;@4<�2on��4+����A12�2�.H�b�����M�������]m�զ�ዘ�0�G��P�@��"�SŚS�_���'��z�{Ǡ�hf�E�,��P�ʚ`@�I#b�c�G����i�ղR�������D�6bITݽY�-������a�A&t��VN�O�]Cu���#��;ZSSZ$�"^<\���	�&VD��9�ag��5�	��t�.��񁨫�dR�h]Ӛ�\��+�@JOhjH�v����/:\�G��s���O���O��8�^*�B�n ���u�3�U���i�B-��nΧ���=���g���c\�@R`�w8���r����da\G/2Ke�rYd�Ť#1���t�l�vR�6��.D�>��D�Uwg����N[Y4��r�4�,i��?�2��2����£��-whG'z���c�*7��T�Jq[܎=̀��^=��8�l��0F������}:�{)\\	�Uk*�D�z6ÛRs@y��b�)�7׃�c=얤8� �X�"�5��1��g��~��C}���K23S������c(��E#0�/���a���&��W\�~T&�L���mm����k��뼀���5�x��a������u��E�j�D��3<O�4Ϻ�eґ�IXB�C_-�RK�nLBEO$Vn�tR���c鋋�5��l%"���Iq���`m�ʛߣ7��θj?'����0���X;�%}(u{�љ<{ͼ�}��}�[��;��"@��m,<�<mc�4�E�su�Q����J0�2鋰e(����ІAb^���7��ţך��W�� :XǍ*��1�a��	�7���
h�!a��_Q�"��}���~�]����PM�=WCP�H��onI#�= P��&����7��QL��2����i:M�f�L�lú8�VK�o�.H��Ya��bKA�F#ʝ���@ߠ7 �
�aM��e����o�kY��(	QzC�+����L�<�+@�xA��L����^Q�jB����1���U�	ߑ��"
�ׁh*��w��gog�&V�$K�zr愖�F��E;b�h܄��K}0�}�����&���dҧ��iw����"2�"��q�0�]�X��и�tw�d6��*A+�W��LP�$�c���Z��;��0�^��Ǝ��_|f#L�����D1�h�0Z������tӃ�ec�H��d���)��3ʝTi ��	��l�7Q%�	^x��o�_�}�FT�6?py6�>1ō.#�h!x��������75�3�Ae�!�ܗ?a�n��D�bw��o���L����f��N!Ү���+rH�j�'9��d��ȥ��ܚ|����:lN�����3��W9�$WYK�0��V-t�\ �uR��-#�	���[�^Ofg/�����R{MԠ����|me�v�{a�垆��;��>M�pP�	u���c)��B�,Tyi�u�����oq7nϴaGި��me�ٔ7�T��_ޒɤG�1���2�},� �7j��}>,7R���5�����GI\��[SD�۩����d�r��D��?�n�H����[����5��"5��J����]�5���>R��I4%�)yq�o��M�bd��E(�f(s��L"Ļ����VH��7-�
�%�-M�8B�X��3:�ɲ���e5��FUC7�+���"m���j�[��c����ٽ��ݏj�����[���G�/4�M�ǵp��P���Iݽ�b,�(�-�@S/|w�������O���� &&�Z�_tشUM\J��5�~4=P�7x@���T5�	&.�{_(�ݢ��Z�[1,J�)!���-#���l��*�Y�J�F�m���	Ϛ�M}˕~���T��Ԇ1�K�a<��l�f�F�c[�aĸ�6�t�_ ���U�g�8���N����/�+Vc�T�r)��ɝ�^�d�p�||
n�4���������[Ŏƙ	^_8�
�r�[�x��R<��)pj�P��-��r�q��̢�G�X3����4'��Wۯq��#|�S��������K��������SA�!��DP��2,��D���$t5�(�ƀ�rks�y~_����@���LkN�F�(˰��#�n�\���0Q��0L}���Yq�2wJ6���xj�`�`??w,p�-S�U������0�����Er�a9����Rk˙�����+�;����q�S��Z������.ĸ�c���:���;�n��\����6<0/<L<I68�D���ڹYz�J5$�֐�	�R�e����(cR�G�-
�Xa��(6SԸl-�[8�jO\��)��dWB�N_�U����s9h���巟P�X���`��z$KJ:�R���zE�'u��z;�������t|X�:��ñ�����s�q��{Ek�r#���F��<�ܜe�L��/CF>%����Q ����>�aZX����O@��ki���~��H�?�)R���BOVC��9y.&���Z��>F�F���[��Z^^�H�g��C?�%��w��_�t���G{4m���q��k!mw˹���������k�2%I8o��2iVE�]�)�@)NT�=w�%�?���X�Q�6�B�Ssg����x6�~K	�����N����2A&&`vU�	����J:���v;h;��I,]��)��@Շ8��a���������6����ϰ!�0,����0߻���v�)��Z�2 �w4���F���=vZ9����Ƴ��t��ƳC��+5�ʼ�Zt��Lr[��{y�QӮ@�⏹vV�X����l�P����&E5�F�\z�|R��i�����&�ʣ$��T��;�M�P�X��,Qy�1#�d�&[�t�߬���������4���#"@�`kez	͔��lChD<�c�����w�XH���..�A
��+d?�L�p^�b|r����\�����)�k~���n7���/�J0'�� ����š��YZ'�c�n�W{Y��r
F�"3+��1ٵ���L�X��U�*���؉*�R��+:,��W�x�k��S���QTG|�od�=\=�W:[;S5 �A���wPl@>���D#�3Z�13��Y��I�l���7P��,M��C��,&�x�d�A��VGH`+&g���y����t��/Q�C�����i��,fW ��	pT��v��\�z�ðV��
7-�j�A���
�;z�.#���5u�l!��jIZ��pذ��v$�n ��Ǳ��@��g�V =�cqdvw�EF�F @oBt-R��xp.zK:0�_	h�Xo �ˠ����ئ���om�r���gݞ���+2���p	�Ђ���l!�l�(��_���|������Z�5>(�(rj�7��A��B;(��`�k=pk'n�%8�,
��o�������_l9J�d�����.�c�����} ���׬��;���$d1�`*�g�x��+�S�>�$7&��t{�͐p��i��� }����i������LF;�;d���q����pR
���垆V��ѩ�Q(J�>���R��{�kLd����^� Wdj�����-*��Ќ@8v���rUQ����~�`� 1Cj��AOI�s���zt�}͕+��������R�I��o��B�.�5�B ��|�,a����ߊ;#��{�3^Vh.w�oT����5��4^���4�dL0�r4����&��'m��塃�3�7�Jf�X�]���f�0<,T��:)_؂�-�g�P��3��l;�6gI�K)�T	J�F]-�hM
�dR���g�V��`'��|����tۡI�36ۣ�"O�ۓiϲ���VG��8Q�᣷F�?���f8y� ,d�J9�福���`�2�(�|r[!��0��/���E�(�#b���χ$�=?�V��:l|�"�ɧ�^h�?�L�B�:Y�X�f��<�Gs�cB�{�ǎ_��7w�`=��F� �B�rf�V�'�S/�P�z����L�?�.C!4L�2ny#G�vI��0�4Y��X<�rKí1%�/-��5�o��|#�.@�	<���:��X�us��8�9l�2�B���{O��f+�\�$u���h�L��b��F�j26�i�,�:����B`��&O��yq�_IPS�q���(^j�e�T�߶�J�Z����ژV�*�o��M�]z�Y�CX���Iq9<�aZ?AN �s�B_�Q�GH�BEp��C��]�@�AC(�n���}�A4�_�_���Bw]��+'���[� �.�PEHBȧ�B=��c"$j���YK�D��>(��# ?6L���4��%�����n&[usm���En\��f���e��pK^���_.�}��х��uɫ�ْDq���*�*C�l��X�]����"�����n���ؿ��"���;Lb'�Ok��<�<��/���(0Mv�m!��33@���,��ϼ��f��?%�o�B��4�0��蝕�ŹG���H��"�{B�Onهg9n�K�� S8(`����x��F�����i=BL�fƍ�������YgMXA��ᡬRG��
k�B��w�>�[��=�7l�U���.���@4舊)�Y+�9�㞉��޹���-��胘<B�b���">����tjD�W�3O�'�_�U6�+�F�V����W�Z��nH�ID�w7N��~:N�}��T-���εT����I�E�/oE�$�����[��_���`B�<怉�uB*�̣}!�rg|�k�a]���+0���3�w��"M;g�����(��2`KD�H+�Z���降��uYZ�Zt���e�YEQ>�S� �k�!TEm���#�HL&�U��"��=슝��Ʌ��~|����څݱ�5�Oet�8/9�#X� �6�"[r�jX�ĸ��%fG��'R�����=x�օӐ����Ԫ�<)4����ľ��W���A!��\&F����ܑ���E�� "�o��z- `���3`��I*��蕱[IK�ոV��T��*��jq�x� q��u�6ܵo���1���è�R�2E�]q?�W�El�]�k��~���+D���(�u�Þٜ�҂KA�J������I^�s9�/v(b��ʖK�#��"�~�Fex&K���Qh���@+hR�duh����� �M�$�R�C�	h8�Z�a��4Q)�e�[`��
T����bH3h�!ZB��B�l�eon��Q�r�����a/�x�:�:!�Fx$b.������F���>z.��/@����f;b�}�Ȅ�f�����,���e_�y�P��*���s"��[t�i�.�����zJ�'͘�4?��)��Q�CD��t~غl*�"�d��߅ک|@�G*��C��`�Z��d�0ʏ�II�M�t�:��nӏ��V��D�b�z�HQ�D+i�@-�C/�-4��yJ�N���B#\�����n�4���=��l_q �;����\�hz����EwI�y"�����-��l�T��|Խ�.�.���>��	F{��:
�`�	�D����c}�ˣ�/�o�hE��� ��)�?7�1E�#9��x�,2����hg�MMPp��bU��A_L��>�.Kx�^���Nn�PZU&zF)$�M�$&�>�٫��~ᲀ]�X����RP��U�GNG����	|K�bJZk@��dS�{��-��v�@}�a�9��Iَp8���a�}�wC�6L���}�L$؁�sFd�1#��쬿l楈h���ÒaF��Y�e�O����}B}�#���)�W���Ɨ�'Ng�jgR����E2Ek��L����H:?�H@>���M
5&ޅH�{�K(i>�Fr%�w�DR�y���K5ߐ�#KݖM����b������7O]\$���}ɿ�	�cըٷ
�Ĩ����� t��s��֔L]��j%�\�*�z9B�)�8�y��,4_�-7C��px��� �
M�=A���w��W|�8���8����	�oH���F:`��o\�a�U�h;Z��+^l�	X����4���Q0٢�5Dw��Mv��`�w��S�u����pUW?7�ף]T����B��HK�n�V
Q@����)|�nf��z{��޸�Z���D�R/t�~38P��bZ����&YX�C�r�qi�,-�7� ��4>u�oWy��@=�0��r�I�8���XȔQw��ް��oS	�"ƤGx��g5���!!���z�nm�^$B-��-T���́#���[J�;F��Ɉ:�h̭�=�"�H�3021�C;�D6Dk�e���5����M(�1Ԟl׾� �Z��e��)y^����*r���r>>1�3&����#�|�P�A�(����"3�63�4�A�lU�����mJ:���Kj�U�n��le�����҇x�kn���qR@�*��9ƈ����<q5c��w�w�c�����M���,xu�lt����Yw����FK���W�Pg|��-�2\d6����GK����ɺ����T��^B>�,Ӷݍ�B/}��W�?����2{�6|&�=�y�XQ����!��&,��ˀ��R��6:#��n� Ǹ���п�G}���o �\��!a�J�I"�"I���؇�v�F�ѥ��u�j��^�f�����,��VBl^��Yc�#⢀f��A�<�=�	�a�-Y�T���Z$:&=%[Ƣ��Bgc�S��X+�e�2�x��P�xm�fs���O�k�?��/��Qۣ�bw}�F�V1�M�1�6�<�'�t "�r�)q�\+����Ib!*K1�\��{��=ǜ��;�p?��ءnګ��*���LC(��/�}G�uT��1OvH� ��آ�U_0)¼G��T"�y�p5���u-���U$P�������_�~���Mҫ�b�֯�"��?��$2=���x�����3��S��wMON�-�*��̊�����=�(8[�0���m��EZ-��@�]�!%S��O� �G.���M�ze)�r�$�@���掚]�9�,��i=�y��I��&����Y�K�����Q�bhӨ���ٍ��M ��i�Y<>�n�5�G�p����������H;�~o��+^�I��QV�~��V��l(O� �O��xJ�[���gWyҸ��Һ�j������`cQC/��#�&�eAA�%�b���[kD^�фc�E�t�Lv�H=��r: �jpf�N�Y4�!����y���=��g
iM��PE�SY�y��j����!�������<H��J9�i�����^E���z��>��Ǎ��6d%<� �!�3�/#�5<y�c!�?�߱�.�{�F�p��y�k߽�]EJ⸹pn����	V$��Yx�������۴�3�/Ym�\c/�8�""�m�%S�L�M�W��Q�P��� �ˊ�E��᯿G�@�-,�X+�O�Z'���W^�)��nfPW[�� 1�#��$��$����=���'V��9��yd�E��\Q����I��!*��*��^-����5��ʆ�
4��S��R� 2�B�kD;Xec���ht�� (B�.5r,>9�D#Q`bt�|�$ip��q��*[��=����/��U�F$p ��ϙ�x�=�^3����(������oY'Ȩ��V�f�S"=tB9X�U
,�x�FG�����fQT�V&괖s�����O�l�����؃�G�O
 
��G���'>-|&����[ʌ�NA��6�h���h��1���]缣<|X��x�ʙL]c�$�t���}�R;Q*C���`�Q��6�zE���o�
v��?��T����4�>�{�!��zӍ� 1J�B6pbu�u/�xRk��K�!� gU���k�;~ۇ��!D��]S�TF�Y�~*��>��A��b�%�>/�����C�e���5��C�q�3/.��a8R�[k7D;ԅף+�,�Z����2H(f1�R���W7�f�?�pG��u~�l?�_���;��Z�a]I�;$9u4B�����a$A<.3Fn��^�lv0v;�zǮ׉��tj���Ո�QI�`��f��kԣ�ig}����{zx�v�[z����T�YL�2��dNg��O���0t�͏�j�'H�鱲k.�hѶ��;�.&������R��wY�>x���BÞ�Bc�Zi�ev�e��y��_4.=ހ�e<zs;�)Hk,��8��D�~4<�(}�o�;��pb/ӑ��2S��Jm���9�T:R�2�p�K��|���+}���m��@ ��*��S�I�����B�
��m�r�u^v�7���M\�H�넧��LV�5�/!�빜6�?Jt:��ly��vI!p�QFg0�X���7,�M��[���'	�k�Φ��ٚ��\�)�l`�(Ԝ5��� �v{Ǉ��E$<�K�C@�h��U�_М�K_J�j�T�V�4_?*V�r��Kʸ-�0ð�L���G��#��_e�p)�=&�7�P�^�j<_�nܨH(vja�ISY�X�@��xEv��%���8e��j�F���#D����F�ԙ��yԲ����D�5�U����~��]���ٹ�
E~�/���uQQ�2J�]���4'���$������Ԩ5�J��z�,��|��Ï���a^�aNQl3Sat~�q��0
�5p�Y2�����ܔ�CA�Be+����9T�YT#gQ0ܨ(�]�W<���>@�[� K���s`z��o֤�lڰM����z �m�|�1�Tf��&e=b��A� 7��Vo�+�(�� ���w cA�ЃᔢXM�S�6v��\5��u�[:��9�?�PxY������w�F�b;­�D�I���?���X�f"�i�����q�HxJ�����¾3<7�̠�� ���u�^
l!���tݝ�.U��譌�a��j
y�tt�F�YBii���ǵ�!wT������:xm���ISq9��M$ʓܱ}rV�A��%��o�x�Fz�͸9 >ٓ�Fx!�[��e��E��������m��ʅ��N�����6?�ST	8�|���B?���65�+nH��'�N�K�[1�n؝��5�to8�%�~���$PV _uU���T��9}��dN�]K�|�D��-N�8_�����C�?�ԌfE�*pM!�a$)�5�ȇ}}����7�u�Ի��t��+%6{D5��[�����6 �`�4F��cH΢��t��/�Lk˒r��c��f�dI��L�b9����k%�]�/�&i�0q�)4��R/Y`�4�~)C^/�>��,&k�\m�m~�+7:P!3����f�������S$�)�@���dP����A_7�˲j �B�i���:�WJ��xUU�U����vGF6��h)�I��d��T�]�+��߸�}��&�#�tM҇�J���&L��P1��C�M�7�~��z�����ԩ)w 
�2?�Vql Ռ-bi/��*�ι}���{G�1�=t����m���0�U4�*N�;�D�*���:I�"�z5VD(��F�j�~�N��iaV][�,h����:�֟���k=�8�ܬoE0��K���o[���0�\1� 9Q&G���λz���a��N5@mY���ʼ|��B�M�-A�t��,g3gU��
F�4���khD'��*18�1A����<�
�-.Qt|�8a)
��;d/����qF�o�l��)	�{��q���
�˔'��j��Hj��G?-�$�;k`U!�7w��Bv�2��Myy���D���m��Vw��9���lH�;�1�*�>���	n��lU������.'�蠙��b�̐_%�$�F��D����*��4��ήS蒝��h��r�Q^�$D��Ns�t���}3��Қ@n� ��ېy�c�]�y�,Xɜ�u��|��C���y��:��P��1\��4�|'�j}m�&�;|��Mf��۶����{i��fpR��F	�<E�����[�>*'�;a�ҿ4o����(��<?�^�L��5yZ�sr���q�����/�W��5�u��:�x���U�ڙ�$;�7kG���������F Hl����3E��1�U�׽���1z^�8�u&��S����GV�=�=9�a��E�v��"��!��@2m�����0����Y��p#��B��	���%d��S�/�F\�Nka��XbF��F�MM��� Yl��K��<�xe�@�K�r��kV�PvF�N�)���6+��<`���yח�C��~�n���f��<MS7$&(��|u���?s8!J����i��}�*K��@��e����u*�!�/4K��O����t��͑�!�ǿh�9��c�ӑ3jj4���xQJ����8�x�E��w���6���r��)B@@~��)�(�Ya�G�ΛܛX7!�6�%(pl��:4]]��iW��\ބm��jeA�>�HX�9��{`��@����0�9�G�-�v��p%�@��[,����GdP;f��9_r�u��S�D��@�E2g�Sh�O���w7�Y�2��Wy�D��d0�,���p[������N�ZMcNT!�"ߒ�.p,�.c�|K�/0�����N�6k$��ye�н|�1�-0$rhw�f~��ÜdŨ?��sWIV��ʁ�ya�$���طrv��5J>�.�V�B)i��4��O8 E��Z��w*�A���ӽGv)Ö�
���$�}fHq��s��\(H����KwX >��oh]k˔�
�?�Ң�%�d	m�\B9����)�H�!�ْ�X��4�xl�rRz滥��R������gk%V!�V�oՏ�t���n]�_`Q��� ����j��I�!�7y%WF����t��L���Oh3���dx=�v�q0�^��4�ÉVo�)�"S�h؊���a0	
P�7�<U������c�"{M<�b���l�0>���J�f,���YA.^?�j���Nڨ4`� w�F(6M�����J}��4<��>�^5��;�̀"Hy�CiH�������ˬ�o)�7�}�A�<��DX����&!����l=��������b���`.����El9���G6��EH�R�z������E&^Y��'^��3l�`'�%�kk���קTl1b� H�ai'�� ����w}Xa�����ng=�Tš��%��8�O�{���FT~�{�_�p��i�����;�~א�J�)��8[4I�!�;R{��0.���1�گm��jt����# r��U%4q�m6E��0?�l������k�����}w.v���L��:P_���
*���%�a��* 6s�x�|����:T�X �V���d��{���6z/Q���5ʙ�)�:��O%"��Ť���*��:�)
E�O\3���O}��O2�k5u�m�G������(�mY�����~�X�o�[�ho0�:9�Qb8v��2�j?��A�P1$�pZ�6Q���P7����ZO�-�xsj��o>�kkp���PV5EZ<���j��{���f�o*���S_+��?�y���!�dČ �o;�bܷ��	��rv�3��������&����K�:�|�Сeo� �����r�:����}�6�&#�W���Am#/�GȰ�n��ong��]��*��@;��Wu�|O�~k�$V$��x-����xE1�Pr1wZ]��������d|z�_�U�ax@g.��B���8Tm�#��g��sE�\S#n������I^���ǅFat.�]�B,� k�MB6�]Dv��&���16����]�Nm�mN43�dAn�� )�uZ�sR~Y˵�����i�Sƃ�b,�S}@M��֬����$��N��,�A��R�sY���I�&
K���G-y�\�8ӄ�/<W~ޓ�t����M���&wh��\�z�1L	�׈�7uX��c=�l��CJ�g#@$C�4<X�X�OV5厪q����@��3fK$F���*.x�2�(�����;�k��j��_#@ܼ�-�ԹÜ����Е�)ѣ�~=Q&ʎ�U[�ة�_�lG��Ulޜf]+J��0��9.�1)�PT}���9.����I� V�jm\�۹ �d��M	!o���]�#�9e�r����/�Ōl���s���jƣ�(��T�D�������ic�m;F�Ir͗�r-2��}a� �ʢ�?���X��'�v|��	W��'4yr&�e��z�,�kk��`����j��(�%����ڣlx�k��K׀̆T/�(!X����3!EmGR�>�F۞����%"�y�����4I�l90)���j�`g����@9O�"�C'E����OTjc���4�$*�#ȿ-!H։;"`��Ɉ!����{B���K9�_�1����7�H�����V)��K� �A�^u�9ސ�h�C��B�"�a�y�6�8:�x�SB(���Ԋn��w/���5�׉S��Kf�rp��+�E�z}�[l��-�Ln��82��Nz FI/�9hB�D�\�ɸ�X�̷��i�<�'��T�,X�}�B�o����FJ�a��c���r���h^��.'�`s�[�q%/XS������A
q���gr�Z�gy�{�Yq��K�ӍC�@0p�}�Fo��/W�ɋ��@t�q���I��/E�h4G�O�C,�
x��_��%B��i{8�q���p�$2�����4���=B
ιbgM��=�K�lJ`�|g,���f�p�;�\�Y�"[V�Ӌ�PP��qV~�!��P�nM�o.υ�o��w����?��\��Rע��|����-t�C���ёa^&l#)��yf��IH���N�#xl��ܚJ����!Pć����<f��[����\�N�E�Q��ն,N}�މI����].�)|�6�(�LӖ����Ex�A]�F��?���f�H�k��SbZ29�S�p�sx<�[��b�M�/:Ne�*<��^��{PR-ELf���#e�xHqs���Yg'��Z�<F�`��±����TMS�O(�EOB pX�E�q9صO~�^{�,=WU�����͝ X�z��q9�����d|���[����z1^���!5�R��Lp��E���췪L��.���13���3�Hx�m��2�m9��V�l�ί��B�Jw�4X!�|*+�JH�p3]yb���)�xM"ѵ�fZ1^�xy��*XN>�3eM�w?�q :�K˓R.�`!֣vp/��!��Q����Ke+MR��y~j�M!�ƴ�Wd��{�N��`ߣ�tc���u"��͘Pm��L��ub��ʐ�Gx1��%�0n%̮�N6v]i�������tc1bX��3d:���0���l� �L9ľu�X_��.�:vO�S�p���n�|��?�,SV�Z_vH]4�NdqF��� �����(Oh�������~�,�W<<��a�,��~��ڕ�-���g�X�In[DR��R��\��	FDH��_Y}�e�7�[��ZBB�a�F�ﳐ�+��R��j^���&�<?�HU;���@k���53}K��u	h	�"��9�
�g31�����G_19���8z��L��/��E����{	�TiWACcV�W��D�D���E������%��UU�<�4�1��\��{����^$� �[P���Ox2�� 0?}��������}b��D���dX �6�z�����?�J�"U�pU�Q��E�k0N�K���r���T����ix!ns�cγ���Y�ʗ�~S�sн2�@�!�`ƻ͘��6�U�/��"��
g��G�}lQU
�G���A��v��K��\���%'n3j:�@v���sm�=��01�I*�In�n`=鸏��HN=,zr�-�<w(K �A���l���a��Ah��� ��o/Y��Ay��)�dU�2������Ѱ�5�;�)� ט��yU�l|�z��	}E�NBߖ밊(�-k�Q�G΃�B�8�����-�Q�ӤIEm���B�{3=n��**4}0���A?t.;%�S0�ꃊ�"	�e�^+*pM��L�e@�Rq��8�L����&7wZJm��A�;g��6�m��t2��ᐴ���״&��?�&�+���yN��g�a\����
��*�'����-�7�2�a����wк�1�5�0g��Ѳ��QG@�b�����<��G��ݟ�O�m�:�����C�Vpd��7ۻ�R�X�O'�U��_�D|�|��yA���r�����ޘ'u�3Aฮ@?�V@�y�yJ���]�5�����Ê��h��T[�t�]���C��Kg�n�����͚�r�,n����s(	Dk-i2���uz�����j�f��h},���ڠŅA�x�����,������C\K���?�I2G�n�1�P�q�;��P�«*v�7�j�M�"<��c�V��ss����s[h{�r�b�,*ho���UY`�Jzz��1#����5|C� �l�k|�WE��k�?��=f;�x��4'�-���G�c�]�"|�^��8o���k��B��W� ���\���Î�;A����y
x`�=��TbӸS�: ��i*)_f�7��і�=�cL??cji��R�c���Hs�vi/_��[������Y�ϩe��B�%��t>Xo��fZ�ǩ�	���B�P�<\�$MB�@e����7ٖQ�{�vL	�)�����9��1��� ��H��ZMK���;�0˩d��p\��;��ĉ��H�<zu�'��R����R����1n��̍��u*�W���*v�~E�Yj����983��IP��m�F�:���x���16 �x����,��DS�$u�̈́}�LkPZu(}v+n;�Z9�,;���*�ΎK�s��� *��[���h��v��{ �V%#���3D?TigN��+{��JF����"��KS�\�)��]�Yq����[�L�?.|Z��M6�R����̡(/���]�S������2��: ��Tt���ϩӈ��B�
�ⱒ���}g-A�4�7a����TڤM rO�:l�OGʰ����d]��ڷ|%C��ʞ��A��\�d�>����uZ�
��r1ڏ����B1���W�He����
g���ԕ����2;c�.q.���ژγ���ޓ��ve���-?��Z� �5�FyH^Y3G�H��wI�`��0s��]��| ��`ۖ��gl,�����o�3B/�gY��a9����!�W�[i?b_���ҔI�&�TP�u��U���+2�bB�52� |�������|�x�7y���G�-!��eh��B}����Ej�����<��*\^GUU�N�c"�"*Գ�9 ��"����@�<�$����}�	��c|Q���2n
W����(��L��L͝�>%�_��79���M�"=��1��j����m�>�.5)䎟�t8�t�>_o�j9�=�D���7���g�}>�U���=��i�1�vhl�~�8=�<�Z�����GP�R9��<�l4���A��'��]�1Hy*0�1�:u&j��i���C��y%:�[v蛈��n+��"w<��Y������h�Kkb�E�9*6�F?$`usA��qw6p6���������q��dV	ēB���|&�9w����QX���g�xG�t8P+Щj.�~�N�S!�Ъ�@͖a1�Ι���~���^'�]�m�n��=P�$���{%�H�]A_��ʜ�-q��m?GG�vm�X`c0��e�z�y�\8�H�'���0�gY���y�� ر��R)�}(��=81�P����d�۬��A��gJ��=%#�XA�M��z,.қw���&�����oGֆ
�f��B\�Km���G�Tg�Ta��`�
c�%�2�|;��8�yz܈4����B���B�낏��l�Sh�?�mY?�'yM�С�s"����/�˖�|�^d��,���7�jz��:v� 1]n�$����_��#��Ɖ[�ɳG֟45��>ږg�q3`��S�_Fv���̎.�������ߏuV!�׿."�s81�J��#Q3�m%�U���e^���`i��@"����1HB����tӾu� ����w�2u�t�\�M6/Gazh�.+So���U�!G��/2�-��q5��7{��J4"7�� G�ZRCI����ϏލE���
��BTY��I��=$ �nzY���@�K����їm3EG���m��&��i�g	=#'���'�$ӊ��H�0� �#6{Q;"Тh��L�����@��v�% i�*.!S��q4 U�@���A8ڌYf ]듙Y^p^�T�Ȱ',c��H҃�,�&+�I�y��>�1^@�w���yν�;.����(��o"���y����W��[h=�f?��3�^E�$#�@���7�kt���pʗ���RG���Wv��әD9��Hi4�e�,���!#F��0��O?������U��߅)�2�ڋ���ǩ�lic������EL�>��b�M��:�2?x��ޭ��l�t�����T*�O9Q����a��eʠb���T�5��i) �S�(�q�����>��tj3z�9b��2t9�x�N�,U�:�(�ׁ��p`�&.�/���!��6m.��^���1b�l���$땀���{N����U}P��ӡ�����ȊF�)���0d���~����e�BTG���t@�Nr�Q�w�8�%���
lCx��]ê��L_�Cߨ�eh0����ڠ<���C��,�q6xu�w�T&�b�p/������ zk��x���2q~�Qv�tk�4��IwWit|���PF�2��j'H�5+�ω �ZW���Zߟ����b��`};z�p�hF�g=�ހ IO�u��w�H�NXV���؋�	I�"��[u�0�`��87� q82Z�+6�/�EȤ�c���kJ���'����Ũ���Sаu>S���q� )`1���*�����U�u�*'�=�0Fɑ���֧ޒ�ŝ�A�4�b���tڈ���S������V�n&�4��ߥ��O:習��O��X#�G�ԹÞp�3,'�n+u��6!���-�ӎD�.���.5A�X��K�V$���.vvS��#��[�먆g�|�7Mo|9���W�5���O+��B��>dbZ���glg��m�yI�͖�ܔw��T\	S��� =���ck�!�X	g���GG�7ti�7ӅV���?³(����{X	x�闵��z> �{(èD_�$�Ҕ���I���F��\�J��zG���tS;S
��q>C�Ω�ؕ�x��rx����x&���>�'�ec��$�3��o��d
�Q~�t�'8,Y�.��.��1ց��Sn��i5�Op��� �"����	M/�]1�:D�� (
]�+Qi������GdRaѽ�M[Ļ���)�	����?i�g�����i��r��B̷�BP�|���{�Z�>��S��x�<�}���bڻR�}1�G#�lxl{�N�yYO���1W�(��,e�~Ra���?�,Y*ɆgJ�$x)sex��qw;J)���f
�����a�	�1�'.�-ߦ�>�&s\� �SN���!y��l_�NՎ,���-�7�/{�����]�I��%�C <��"�|�ݍV�Y��Ts<��D2Cwfnޡ�l�Dn>&ʺ/n�?�t�(�d��T��	��Z��X�&=$��$j�� ��Y�������?S1NG��=+��AV���>� �MΈ'\az<n[��pq�Z��B��U������Ȯ�L�K�ǪC�ۮ�Pಐ�*��eǏ�s�����{��LH�̰u179�]�8<3d9�?�����C�������F��SF����l;N���2M�V48T?�M�y�����6���t��b��cIF<t�xS�p�6�R�^�@6[<=2M���C�̌��F�u�\�BK_ݽd�|2X���htNL@���~mA�=Q�V~�_�뼱{�C��Ն�����'C���(1�>��]=��%t_��I��P�'��y���w��s�#���	f�|�� �~	Cn+���]��l�Ls�6�^��kJ������b�Z e׽ԅ���N�p�3�#)��!Ac �kϖ/Q=u�
پ����m�\�#n�.�U�M����ȼ���l�6�M�:�E�G��Wu�pV������:	1�pT%
�*N����{H@���Ka-x��pP4� ��`m�����A�H�$��-gB��PZy��-�o�1T��ku2(q����ƒ�κ��@P����P*j�0�F�_d�86 e�9�����ߔ8���u������I�/���;�����(=��Ou�T�����{�ڃ(���ݚ���s�@��.��eQ2��q�V�U�.j��������"H��w��,�vf�or�!�]Ha��v���f�:}��j>*�c��u:?��O��7�.i���.�|�%��$�	�q���L����4�?
J�ѽ��h{�aM��ѐ���$p��K8���99[�G��I��^YL�7����N��x����{u0�JS7Me=Q�{f�E����a� ��֧&�w)В�Es�Q�u�
&�O�ao�=�#_�Y�м-�� �
�V��lF�5�ֽ#=@q$ܕ���)/����,�S�=�\��mh���_�~�S7Y|;o�|�M�\�p	Y^}P���$��e��9��b��{J��dl�o7��׻7}���P���X����eiZ�Y��K(��@> !��.���X���BK��'TYB�������I%l]��h׈AՆx�ӳ9:uC�өh���T:@�,(:�v`�?�(*t�-um�=�M��M��ޑS�w�X%�l��^��X4��!s�Zʮ��DF��m>�Y��q'�`!�a�>�j�:���?Q��@�,H�b��\ol�b���\qu2�Ϳ8[0������^��2!��&pf�]@p��*$��
Q�]aw���GoQwX�������h>��s�F�K����oH]�[�6��?�9�0����b�oz�2ܻ6�q%�eє3����Va��R<=�0�0o:��W����b���|��{h��+�DT���
�@ց-��P���n�@�����7��K��[�����'t����R�2e���W�s̟O�?U��jʆvi>��SG�sA良pxྕ�ۊQ��\C��c��oฉ�
�ռ׍!1�ͪ�{ȼ��"H����#`��&5+L���K+�kmv0�l��@��(i��`ȃr?��n8h[#Ň�%����QX��c��=�A���TMŏ0HѪh�	m�@|��$��lt�'�*,=Q��Xʟ�*����f�q�~�$*6���ۅ���7z'�cm';Q:`t���\�4�:<����&p�0;TG�H����*蜯�R�S��AkN14��#�읾Aŕ���|�\�Ji���2t��_.�o���
�e�D��R?@����\ ��"���0�t���	�u�֜qS(L�f8i�K�E��w,]�]p�d��'[�����y&nY.�1�;`l �62Գ	0�2�C�b|X���J�T�BVI�p�Oh�2w��x]�(���� ~*�����<2�,�#��u��&���}�2G��/��X-�e�MF�� 7������7�e]	�.��; ���d�Ĺ�-ù�� ܪ+"�L�Qξp��f���t��_p�N��`�e�h����yj9�K<�p��� C����&	�@K�a���Te�7꽐��8 u�pD��t�gQ�����RQ;^�uL�!a���W�r�q|���LXUI��5�wA�5 �W��,|��NK~�u�9��������1Ŀk_`�ek�P����g4=�0�����R��H�${�%���x�Ï[�Y�^�v#O=D�dS�h+��xx5A1B�4�����uَ�$�����9�!���ꄡ�T��*]�@�P&�j[���{�t��G�Z��T]��g�F�{мC�	�Zؓ7�q�����f�;V��	���%�^�}�q2�D-Z����
�[�nv�&"/d�|��cj�{�|�v�H��Uq�Uڴ�X�X/ۋ���HE�yV�JVuT�������1I��������Ư�E�_���x9�[:�)�d�ŀ���!I8u�qJ���nUAv�F��Tkꈵ��@�N%5/w��ڭ~�C'���|����o��R7���'uKC��5�L�TT�2m.�Qk���:w���*5dM2.u�FK8��;�|I�܄7�G
[��]8�B2G���q}b��Uy�>"@�����L4@�?Āy��׶;)��Utԍ��I�vMa=	�%���`�וP3�,%z�@��~\�JT�惩m;����fFs'Ѿ�$L��u�]����惵,@�m�%�_���nհ36�d���cvd�~ݩZ�yi׽��cP~�Q�u�[Em��PG�W�]x��"�n�s7���d����X�=I��eD�(�pf' ���htq����p����K�b�.��9�]�\ �(qZ�v��C��ZMk�P~�Yޠʛt��m�ǻ� #�\XY�U���-�#���sJ'�,���A�|2����}�cm�T�)p��@yQ� Ï�"g`�Z��@.!�,���n��y���j�9��#����#8�)xc.{^�H�d5��[��]yӤz��k��۫#}�ȫ;�DD�u���s�%#���^�n���Yr%ڽR[���a�j�(�X|_+��d��7�aV�˭�����^�ӫ_#"�
�o�\`���KO���8�8¶��eA�zڣa�N1({s$�iL���A;아���ϥ�t���x��liN6�k��e�ͽ,@b 
�s)o ����rh��B�:Ӓ� *)�I��G+����ܒ��k��O�3XS��3
$��)���c��o}��`��m�*q�[��2�J�~/����K� ��#�rVY$}�uq�
;����Q�>=�!芢/��TMN]̢�&��%y�� RRf�����0�{����J�\N+<���⣸�I��8��]���a���U�6]�M�۵����"���i1:Q����ؗY`Qۤ�P��e����;�[��#�J��yȘ�߈6Q�f�=5��՘�E�}�h�+����` /w���h��0je#4ռ�ƔS�)��ٹH�C*�d=pÌ�E	'��_��.�53����;��=(I9�:K��8�8�/��n��dhN&�����I)p�*���8����:|��F� e��:>��@�# M�p"BH �ý�D�#�H�-�]����$2�t�:l]&�D��$Ɖ�F�Y]ch��.Q���W�0\�^�|LUV����t�ù�R�ߕ�TԧS�����F,ɋe�E 3�����c��.��[+W|8����:6Mu�8� ���!���7���1�9
g6&��vo05�	��J�g���3�����r��8�s�B���%��
ZI��H���-E9���]�))5�v���!��c�����_A��Jg�~�'j���1�|��M�V���l3��$m�m��j�Xe���/c��EcT'�zӟyd���dl��y|��YL����J����������-�֫��z�xƼ{ZU2�xd���{^�����{�����|
��x�<{�]i�:��9��Z������3"P�o{�9����D�s�?VX�����a�W�zl�qD�w�����\<���Q_a��9l�a1�f0H�8��\bp�a��_Ƴd��C=��F��&+ �t���0�t뤟-^�7x>n��Sor��Q�p���~���������B�F�`�����4��V�4Ϋ˵z���-����&3��<��Lt�4C�{���VR�'0V��#�����?���]uR�-�=,R�K!������/$Y�����٦����hgj4Q�$�wH����"D"y�Z)�i�ގ :�����Γۛ�Q��C7H,��O�˽hOw��?X���� ��eΔ��ݐ;�.�t��u�ʘLM�W&+���zI�ޜY��yIv�'�L�'C���ϸ;`�Jœڣ|��� �����ï��0<A(���ҋ�u�fW����M�Q��d����|��V��g��|,�K��uA��a�H`���s��\�	S�m����h��C0����s��xmi+�i��Ԙ���)�DE伵��©�S��]���S����/�@e�=�Eez8�?K������.��AT%�3�MḠ�o�u;p� ��8� <��z2�n�Ϣ�)îO���W ���ǠW�����K� ��w�H%@��zP ?T�xUt�c���ayH���W�k�̾>^��.e��Em3߸��X����ַ�^�f�]��>ù蕄B9�	�}<��M�M��;ߴф��?�Z�[ʢu �H��T���.�>{rg��[,ü���,0Թ��N�f���`��a�R��8�4˶�3<�&�ܗ�T �:�<hСDO(j��Gg��DD˕�ݡ �WR����q�l)ĺj����K�Y�������Qj��k��&6��I�ZO>d�m��7�=Z��a)�+e�r!Դ�X�7e� �GӶܤ���Q�κ�mIQeAW�!��DJ��$����1de^�e$/�fs'�_~B�(m�F�^	)D������ǭY�,��p[F��ػ���G���@dV�в&=WV�����o{2�m6���J�qJl��fI����u�!x��G�@0m����RMO��o��@,�M`�Gj����GuO���=n7
ǔi��! ��Cb��Ċ ���4�px*�7�蚉\���0������H����ѷ���ʗ6FN("(oC HW6�˪M5��?D����^��ItC짹g�d�tp6t�Z1Z`��͸gݼH������	bi}�R��U�����4��R��"�Ie�:�Gp�`�{)ai鬾�y����x�nN������C���NzT]
諴U�
�qSE���[�Ɛ[���ٿB���.B��i��I1E^��~���PnFX�{-gB�ɇ=@f�[4�O����Z��_�%����0峮k,ӭ�$<oIBK����0�Q�Sp�$�f>��������v훥�zb`�����)"\�#%YB��2�9@�i?��r$��\��T�lq�%�G~|���ɢCKo^����4���AbJ�q�UZ���\�J��]�`d�rs��AY|�Q��T�IO9������A���ђ ��ȟ����5&�ȯ����Dd/?<ѭ�>��@Ӯ��*�lbx��N���Z/�Q��,��Ȩ����
�>j����mў��U� (4΢L�1���h�v:J:�w�b��h�U�*���0��M�ьp��W�i��ͯ��è�$A_��57xp^�	v�J@\�Y���k�Z�u��~"Ó�ƹ�kM-0[����"��̞������H�z-�������K��p�y#}��Fs��ܿ�5��UP�ʟ���Fſ4paRfu@7*�:1N����J �\/��˃����|���)�m���a=8�$���':�V��0�/�X���{��t���JH&�3d����ʷƿ�9�@*��v5&�ӊ�j�F�5!���+~r��
�r�2W�L�ڲ����M`�$M.����x(��" ��o@$��k�:�#=�#�ԙ���H"*�pM��б`F�u����͊�S�,,�؋j	�����:�kj�J׾t��?_աlu��!�#��������T��'L��4�} �^�`��f�Je��47	�c�G
���Vv��&��0���Vy�
�vR�@?�c;+v��hR?#0��m�����[�B�L��5&�n"�/n��Y�?�گ�Aw��wR���@Q��h���.�	`'�jPz��^��
w�,��N�^���+2uΆ�"rXkH@F��M�k��@��4L)�����/��J��;��d�y���c䢗�	�=p�z��;��|O�V���(�铋�,S��\d$��4�J�����}�X�y%i������>m�)��k#��_��z�\�?C��䵠=/�<CAPf�_k��y˓�+sy��kO�5HOޤ�����@l0/�8������P��	���Y4~�~�5�CzOzC�=f�{��NP�+%�Ğ�ە��w�I��[������U?[`�ձ�|1<���U:�ƅ J�V�	�h�֤T�g�jxw�;I#�,�`��@�T�������<fdO�Ԇ�p���p�L�SC��*�\)�DC 5#C����XҐa*����F�P��6,c����>w�\�_��$y�o���-6����ېЛ�~�|�k�!��F�T�%b� 3�4�[��j��/N>D�}V�N)�@<6Z��AO�W�D���P��H�v2�=ʧ_	$ ��I%��b�C���T��<n3��4$���[N����ϤҝЌ+��5��)e�ּz%F"c��T[Zb��F�P��\h(��1��Z�����W@�|����,Ng�1Zϣ2�^�#���a��>k'7=�N=M���"s'�P��L)YP'K�W���篲g(��y!�p��������Ivs;�1����%Tz�z��E.d���l�*���7/��?����%i	3S��O����V0]��UN��Q�>)B?�j=/HIܔ8|�|3Yl揽��cV�E�5\ybz��\�f�5��!���51�.���EPj�C�r[��:$��e�+����\��h�zc�>�Y�,}�C�|DK����}@��k�H���X3�=�ⳝ8V.|�c�b�Z7p���B��X�î�T�s�%\au���hr=X��# \Z�Ls��7tɖ�dL��Y�`Y4������d(���%uJ&��J]����ݶ�w}�%X$z��,�g�b��;���)p������w-g�8�^����,�?��׫_x�@;�>��z�����/�!���F}����5�F�i�YA�^���N��t�Y�51��-#�^6 ǌ��x�K	�欋`09�����5b�\��m�(R�IϥZdy �W��y_�V�S�h�,��:��A`�Vq���4Z��f� i|���Š�w0�?; =�!��վ����{z	���z̦�ͱ#m�t��N�b*���J�H��\#`1:&�ߪv��?�\~�!S	��==�t��
��<�tmw� �K�V0bD��߇m�K ���8��z�]�;G��	�6	B�
1�H��W�bK~Gmv�qր�}��"�ɲ��i���MSDc9'�s���Ӧ���@1��6w�.�xSB�o�}^�Zj��:�VF]�ԣ�1�+V9�¾�AV=���H�O?3��qJ�i-�d$���"b���/�ё��� 9�e,�{\;BݚotW����29�������ψ�.~�$�]�˪Q ��S���N��S�e���ؕ�H鵎Ji�D{�Un�����q�^��UI�>�����I�(�F6��@@�,����qjB�m�i�����p-2_�G�����ڊ��>�)W�_7d9v+D4#�����91����O���N=(�I2�--�`�C�q���}>yH/zS����L�|������Hl�P�ژ�1�n��3дn�	S��pD�Y
�F�r��3�f5��Z�f�2��5�f�|��=��Y��FIl/�vZĠ���X��pNgP��W~�N5�N��uܤ���k|��z�!v�%�2��L�ᇥyWII�|A��u��5�WHe�����򉼭#m�r�Jiy����(�e�*�����6�"�3�w
��Y=h!��ߣ��D]<�9.����Q�������z}�AB�g�iP'-Q#q�+�ۓ���1����� r�BL�����J���3H攩i��JldK�s�2����g����vop�[Z��5�nF�ʙ��o�\�ؐ�v��OT׏����#��/ ��au��b˂Ńs�Ԭ�S�#�lJ��!vA�x+�r�Nku�����Ϸ���?�:���rU�E�L�봞fF�/@��]��TW��ŐX� rZ5�3U#::4���]�&h������7z�LNm�-���$�:4TH����.$ԝpv��L��"td��fķ<K�B�7�+�ݍqj�0��L���ڴ��<}s��:��1B���v�D��'�y^.�ًQ�R& �/��V�-T>�_���*��g��o.��� u�Z��{�ӐyZ�"�����Oq�x�E��=�����ٓ�<1�ض��ӻ����PУ��������nޛ�U���CP�.�0i^�XV'��Q!_��"&@���jEQz�Y|LD���#�8)�@�ئQ[�7��������P���؏�@qO}0�D8|�m^��1)Y^i�����`���ߛ3!TSq+�(�l���]�pT]ܼP$�g~�<R�����*$C�NQ����$�1�R�N}Ϗk�:U��mt��e8��/�ܤV����妨vKt	�; <ꍻdx�ڬ�����/1H�ɶ��kk���s4��T����D����/���҃�?#��H�Yw�NP��7G�5[X�4�b	6�vv%n��fo��}�$�?������b���t�4��/|>v�A /d�{�)�
R1�{��y���ȎW�&u��؊<d$:}9�O�#�T��٘P��7��^�`5t�D:�ۛ}��7@�*z��?�R�m�O3gE^rd�s~��̖Tmt��2X�
^����7���Sg����&AJ��
��֐�倊��SA���KI�ޖ�����ƒ��e�)&������ى`���D�6�61�E��#Uΰ��$:凓�x<�K`D��aZ=��'hc�%NI�E�����V���5 ф�J�ǆ��.cHWP�X�k�m�8�cB*ʬ��� }��Տ�Qﾜ�Yp�tE�0�A�ƭ�d�qp%�$������(/�:�
�zu�@ԑ���L��c3���K�OזK�-�js>s��RI%2ۛaLyCx�tbq�5AsG�B͌�t�vOga��
��pq\���@B��I���F��c$��_ˏ�\�Ŭa��d�n�ݢ�&�ɱ����Yگ��%�r�߅��[���2�v���$7�#V�j� ��d�	�$�3��2���q��e�+ɍ�/�t#�^sT$ff�v��>�~�;pKE��՝?a�ʹRs��Q^��`���X����u3}#{�;�J��4�[]J\`$ݮ�6����L���ri՘f; 'ʊ^�0�� _��׺��ׁj=S������[P�ɯ.���&BM�l�gK���UE���c�3��lߘ�:%��ѣ�S��6�8�l�^(�*�Ϟ|�*9�q#��&���Q��l��_�J�]DA;��;,;�J���@�t5҆�m��}����k��K��N!��7RN�9:#��Mߦ,'\N6ʇ���W�r0{��������oL����1�5T�g�IWb���b���,����h�|���	�I`�-lɂ�--�ɠ�,��o�C6������f�{��:��ќ�(\���W���ӂ���ng��<��d�g�:�EA1�Ky�MrWN<�Ko��,g!<h��Z5j��S�����0˘|�y&9H�C�^���[�WP(-�O��ӕޠ��gG�h��-V�n����r��Ycl!�*¹"uA�	��H�ph��R�je��#�����B򚨦ާe��Zs�7��$q?��i2T׸< �<7�{ڿBΡW ����a<����[ �>m�ƙ��#'T��>�0��A��TQE=s��Д����Iɘf������ѯB�}��s�`}�j�{�K����m��"-���00p95��0i�'!t{�� Ʀ�M�e�ɋ�OCG��5��&(�dĘ�/Wk���5̙�/�uT0�PX�� A	n]hcZ��6�1CM���ϰ��*ZA���w?L1Qs�fF!���WSN"��zs���݇O��1��NyqGP�-�x��Nߠ�It�]�]f���'����'���4X}�@��g����Ŕ~Cm�f4���"ބ�`�{��|��yv�Wa�Ԑ�n-h�H�g�8C�� �]�7/�6<ذ&���۟��,<��
��Dnu�bư.:'�`�\������M���L,՜�`��KB)�H+��㨷>�� W`m5����;Iu?$4O�#> ���q�.58�sF�z砖J6�T,!h"����(2	CۭK 5/��,��}����e&٥�O��d�u�/�N�Q�Ō��ψ^�V��w��;�Svg��/����P{���P���6C���á�Hm>�(]�����B:)������pn��-���.˟�oy(�x��Eg��dJ�{j7�����P�����H�Y��}dy(���a���|��T4�^D�v�yf"��:t�������Vn��g�u#�ƣ��Έ��"$����;`� ��:��y��:{� +Ӝ4��C��YP��e�[7P��n��q���@D���Z�"����d<�.��-P5`�-�;��������҂��N��}G�r%31���|��eB(��03�=�,�c���&Ѫ�5S�繂����h7�"�(j�d�aI{	��ބZ�4*�(�-������Հ���OH�j&;���XZ�u�6�(!��q'n��}��f����`�r�s}�y"�7�hMO�qW2D"���s�J�s�N2ܩ���� 0v�4�F^��|5۽�c��P�x�Bm僈o�k�}��@BF��mRL �2��}!A����s������,�smg8��ҡ�w��re{*�)mm�M���Twxi%tg4X��Y��2�Oµ��n�_�	�Yn"�X��mQ ��Q���a`-��fT�{(ao�T�.�ҬH�w\3��W21�������ߥ����Z���w�ݩVl�l�돈��C�2�w��G�O�s�WW��$L�<��4�O�S��ꕉG�=��N*K��8�\�ι���ޒ--.p��EI�h��!�"����o"���tu����T�'c/m���&v��q�J���nl�;Z�����z��)�t�$i�5D����wF��`?/���c�G�)��yk��>&��*ym1�q=�G��*�~m�6K�\��ޖƠ
p-}�.i�J��B���َ&"���3��SƏ,N,�t9���!!�/��Jd��ƹ��bQ=�'������_��_H�7H�Gī:U��S"`�+�۴�-�w��Eb&�1�Z�6J�De=��8{�������!{/���5>���z�_J	�0k�у@{+y��/�#�c@�۸~���u7�:��DK�bT�%0���bq�Ӫ_��)|�Ѻ���Բ��y;[y,��	(�����{> S��<3�2�
d��ׂ�b,���>%VjAgc�)��e�<6�=:��Ul�i���\Xߔ���!"�p�0U0��Tz�#���Ǥ���FS�J�M��0��RƂP��`����(��y8��w��!�6пl�[(N��^Z\��x2�zJݏ�?��e�2t��-rϊ4sa��6�\����Ǹ�'?������]�xp.�L���Xu�cy��ʊe�WwJ��#=��A/(��������&�:K�P$_�6w����o�'_E��/<^���ӳ��*r ���
�kF�c(�J��r݅[�5������A�4K���0�B�5�/Tʻ�L�Yyi���/�g�0�:mu�SF�4��n��%S�l���)6<�W��h�[�u�_�NJ�e�D\��9pXrel�N�#���Lp��&��Md�B�L���wU��������@t�/|cL���_���0��i�[�O��m���� ��W�ɭT���|Y��U�9J}��J�ش:2�<Btl6�T˅����`�c9L��]Ք���.ñ�9X����Wz�΋JH���$r󀗐��/�R�6Z���C$+���RD6��97��34xc3�~&C��k��=@JLvW��#�j?�2�qDxC	�Ћ6�9{��H�{���U�kU�uJ�ڢ��N @_�t6�����h Tԑ�_�����>��(��st�o}yy�/m����CJsz"(!���d~����Kt�����A��Lc �
�oj���<hުE#������Y����'�G^=e�](�������VJ��s �BLŇ\:�!NO�O�24�쓰��$1�/zÏx��S��1z������c�u���5$w��ǃ�����~w{�d\���}��7��(`�sj������wIu�^M/���m�����E+�K6�2rH�s��t1��A����c�<���F��vȄ��}D���Gr����'l&�W\C�^w6�~����K{BZe�p���Zc^���h��G�DVYf��!�V{�#{�8U�O���������6�@۴Œ�p��A0k�����ʍP��J�L��74wO���x�Q��F>���[���+�������C彴�s�V���rF��#���5L̈́���ym�x)�$=i79��U|)Aԟ�i��O������!y\#~Կtp$21��j��Q�=�W?gyiA%X�W��<��qN���2.��!�:7����(
j{��yʅ"%r���ߙ:�g��P��r�,L���Z6s�_�)�&T��2],)�[>a�(���ڊE ��U�b^���{2DAp�H��jm��vb8�dV ~AS�{=��������*� A�\Հ���6w�.��sE �Jl��넘�J�� ���'h?5ưƨ��_�ğb�W@���W��D�uZ���_��զ�
-��IvƱ�ӹ[og�_�©����]�9�F��hڏ ,�<��t��,]�S|Ɯ|Y�@�˭����^��%����ȑ짅.c�?;�1fU������Kz�h���ims u��TWP(�'��'s���7����:B�������Ż���j�!U��6��KW����ars�����b���Jk��E��i�Q'��F�~������Q".�u4�&ܶ�E*R]���P��^׵>C�*�tmq�V@'8��K:#T�H��Z�Xy�t�ܤ3����f�j�2����kc���Ao�;�ZG��Jj~v�j��)�P��q[&�|�rlsɯ�r}�[���'TJ�����;�RbI�ˮ�}B���I�kHh��b��c�d��aKq�N{�	����3I��|w�شyw��^rn^��`�,\
�V��x��SL¯lG�uv`�hY�fB~?�WLD�Y���c�'Q2���$�ڶ���r��Gs�N��eaQ10��j'�`�?�)��G�`jLO�0�yX��fa����P��a��y���7/���	��6��)��ZBt�	��+�3RlV��\�P��Wܵ,(�]Xڙ"���o��B�������f�(� �Jf�Q���Jx�v�4"�#eH���p'c�R��a��;������8E�;�!K ����٠![���Rj�R��O�/H�����H�Hh���}�����\V`*�.��} �fTíEWD���(f��W�9I��U��zŻ|w�pӰ��}-c�3p�A9`'����7���<Q�p"�<�}�_�4�v9��ɦ�H��%p���2=�H��Ќ��J���:1�k�7yd�!M��������C�&J��5�p�lsMEH=����.���
�)��x��-�R����pe�i^����7l �#��b0Kr��>r���#;�\Le>wˋ�h��ݘ��OK�j��yB�D�*2�d��!��M�F(�۩��U���o�6�̝\��e'gm��5�n�7m��,І^+~��!?��
�|�π��5N%�,;��X�E�Ӧ�"M��u��g
���%-_�O�B\D���Ҵ����%(r�nH՛�I�o���o)]��Z��=�����{���q�K�(ͳh9Ы�a��]� �f�/��} G���%�ͪ�H1��g0��X��S�����^N�	Q�^��Q�Ղ�"%^��+Y�4��<�
�!?�m�r�^����8 ��4��!��'�l�^g�C�緻G���_v�������ٝ�����j\x,��a�8�DL�����]NO~w��M�[���
�����=��+)�wd��Dr��l��z��#�g|�?���Vٍ�&��:qc!��&^�~�&��nD#	tO����N2��PQZ/t**%i�͢~<��6Y="�}p������)S�"kRD�h��.9	Մ#�d���D�i�y�:c?�c��b!�=ܼg��P���-Al�V��M�y��kO�jM�
�ت[�qw(�ڕ�L��%�
s�����2�E|=� ����ãs��Fu='~PftKw��()�v`���fho��:�k�F���'��!02`N�>,���������%��BM��u{����.���"�ǀ�Ր>��Eյ����Uv	~8�����0�Ъ�h}�e�d����psq%f�#敺Nc�ּ!��ь�o��u����k���P���Ƨ��]��L�v9��y_2#�DD��#<Y�C�63�h��PIV��?�*�xD�P��Ö*FZ�z��Q�Z�]� r�@�����	�O�%c��>!!�S����}<���?��|��g���]�Ne�6	8��L�����Kt�r�����V<��O�ykA��Zs ���s��Xe �.�>��gIY=�~�΄�=G@U/��1oIW&=[b�ֹS�5IpD�6~�بC��\�rDfk&���m#�`r�PA'Hi�3�IP�)��g:�	���8���D�fi��Ȉ����^����_W��ީ�]��	��켺@�l�5�"��&k�Ibu���R"5Y�r^y^�>�K��蹃rH-c-+x7�K����v69�8(�6٨M.�6��c�/�4���#���Y������'1}��d�w-�<CѾ�}�a�6#�'��|��}���n�r{�9���M��F�ʌ���{5��5O�v?��.UŃPX����n58��ҡ����Z!��qI�lų�c8��#�����M.<x�x�&�}{rK�5P��6hB���T�ʍ� �<t������������}>6�^��W��(�S����LB(��{���o/s�@o��M������Z�iJu���l��nV�&�/�`��cw�L-�U�ِC���w6�e���]�������~�d��B�íyJ�$}�k�ʖJ?�J2i Q�zDl�����3����cM]��j/;���G���5m�W��Ę��e���Jȱ�����$b��>���`{+Y��� ?|d�;��?��?�>2�t� :�k��2s?;��o��%z�Cǽ#|��ug�F�:���a��d�Zug)���V{��o;)oSs�����Ss�^W��f�@,��v��%��њV�ېǦ(���h�cL[Q�IQr7�4��4��
}8Ə�-�}�f[1�Y����d=�롪��Q�h��a���1J�����J���Yx�_�Aؼn�&�ROm�-F��8�#�p�$
��v��a�΅��}����"�Q���obR�6\�Ue�du�\�2���s���Ek�(w����f�l܉Zp�q_�]ĀpN���6�n����#��p�L�q)�U�]0*6�Vn��`�.1��mq���5Ƨl�LB)���}����gc,-Au^�����"��VZ��?8��6�3��_[P�]����d�瓝�Z��:e���vb[��
�Ө;U�wJ������r�l`(��9z#ُ��m�㧫������wĐ'�u��~bP�	oMÕ�a"QP�`�� y{�5��0̒:BnA�O��?���;�|Z�����x0��QO|V�q��@�&�������i�*J�:�T���tP
�r}�R���~�պA���)�����o}K¾-�}�wY�l9�n�v[6��ی'�4/R�4@�L�J�F'	�<pp�t�A��ԑ;*�~P�K��i_p�خE�CH��l�ɒ�2z�4�/�7!h�RJ �o�HP��o�.��hH�Q�3a���D��4|�;C�,

�?PV`xR�c}�'^Q��GۂJx�w>���6�C�3��wNQF�'���)PE�����K�Ђ�mod������|�����������L��/���%Q5IkYȖ�sŗ�v�ū�����=���W���g��>
8´�� Lc��W'\��H�Ռ4ܜ[�^���'mhlY2P8����q�ۘ�;T����m��|��PN�`	S��K��Q'�|�CչŒ����4	�]3��mj���k�w����������1���'���� �Ǿ��2����R���a|����ZlV�4� �'n�|�ҹ$cPf��#9SN$sه��d4�r�T��׳u��-��!a(-��������%X4�ovlEV�?pf7��G�����@wxa��5~��n+��j��o��Eڜ�z >u�o
{��_̔��9�Q�k�K�-����$�j(8x�\��~��n�X�,�=�-r3p?�1m�r�[42=��R��)Z�C�nJe��Y`Ęև�8X�����x�Ԉ�'b\ �m"���O=�O��D� J,��:4�w������6z��i��C-�S�#�&����
�V��� ��]��)d3��ȓ���L�.Q[,�����g �������%
$�˃j��
mIٳδy(H�w�F��)z�'�Tf�SUt%A^���+�j��$u�H4܀��;��XI��k �R4��ȳ�@����u`��Juxwӛ�2�Q �ӥ0�7 d��	x\����
�����򙣓ʚ`}��6����:zw�6&��l���V��7C�l��j�S!�ɔ����!,��gM�E]3���9Wc|S �{�[�bw�:"�����	i�F��wi��&�|o	��,��t��o� �*�՝���,���	z������=)
�&*��2U�D!*���U�~N����"0P��X����l�Hf��^n�BW1�x��S)�e�
�?oU��a5C4�C蚂O|e���p���ir`��.I~�C����gp��sC�]����9~<Y��+}?�#g�#n���0�w��s�Nώ�, ��.������dޙ�)V���;�Q/`I�j�����j�v3�e$�*�'�Aw����4��� ���
6�Ƥt~+k[L>d���>���$o�]:
�E7rJ�����ɽEv�On����]���VL��mqhS��)��fn[U�Ъ��@w���=w�v����v�V1�P�iB��`���U؀�'�<��yp���p�7�z~�~>>����i����B�m��V��e �b�����Ä�@��D�o��6�.��Q%�X;���y�����W	�4��BN��sXf�E�"R�'i�.� ?	�įl��@'�I�:��AVݝ��i�g}+���9��s���\{బ�w�������Lt	�D.�|+a�킛�b�`U��UM�C��[@��gS��o�8�����J��<�:���܈�βbw3��d�T=���~���Vy��������I�J.��i�2�G����U�L�x�Zݥ���������.hٌP�wrA��I�^����hwxi[�؞���U#Zy�21FY?�x�rK������}�-/^}�*���Ph�h�`M#bg�z�x9�h�s^��	h��7K#�b9���(�D��3x��];9�����k}��M��=�t2r
����c:(�S�44���[�!�A���2��쥛������P�a��T]0���1��i�L����\o���Yl��ȝLd��ص�K��N~�SQ4�Z�բ�Ɗ���F�Dv�:�,���������gvW��S��UW��v�t`�`-t2�~yr�S���8�\Q�~'͚��h[��ny��+6>#�h:�<L��YSϟ��
�����Q�|��A��y����g;���l���[��x�&�q��>`�����5gȘּ��I
�{-z�Y_���T⡸xޱԈ*Q�_Ҿ�i7�dI�]C�]�I$/lJ����$`/g�����h"�E#��9��wW��*yd�E�k��!��l�e�7�� \��u���	G�	��-�[��h�e����C��qq�Ge^,��\���e+�BC6P�c#�dȐ�����ݘ������!��my=t��A��ܯ�hE�N9[�E:��lC���^D1w�p�^H�g��D4��
 �6�ٷ?;�B0�>�[烧]�SE]���ݾ:����k|K��޻B��"��v�(X@��c
*�He�C� �p�<���DBI>�s��}�D��86��5�����h~}�('� ��ë���e�;���&�8|������`��'��9V"�b!�<\�xx!��zۈ8�;���yTz&�k��3�x1���ɴ��z�9�@�� ��3
���5���-r�4�
�m]�'��]H!YB���w.2z����
:c�DS;��c�{E��S��{�jT~f2�̘VɃ���<���(CC����7�Ӟ�~���EM 5�3�x1��H�%���GTb}D�VE0-MF�i;Խ�;��h�ປw(Rټ����MZр��3����eRDR�<ߪ�6���+s�甚rrRQ��#A稰�P�
|5�b�Y\R�t������טּօ�j+x����A9���`�"��9H�l�G���*]e���3�Í>��1�tm��+-���t���xS��m��#�L-����wԧ�Y֛H�M<�,�B��Q�t�ּ�2G�n���ԺWXOzB[�9ȱ��KC��4�Tvx�&؇��������{�*���Q�*��,7���XE�`l��p�΂�!��x��?��P��x�;�q��Z��j&%�׈�G��'+he�Ԁ��Ze3�#4���M�:�Y��"�;P*B�6�n�o�TefB�)�%����$�-�b��yn+D����q�m�95A/��A>B��H�a�{�Q=��
��)��W7l�/���Ru��T`��+ז��.N�7=�K�ꖶ�!w{��(��i�䘧�>�ri��`�hͭ����>H;�D���=��#�ܓ�ö�˵�b�O�0]�g�g/a�gx�����e<��%��+
��O%���GT�&����<��bd7@,�;��T+�g����G��>��If�-	��gf��S�a�����'�j���.�J�y5=$�吶��+�J��)n� �{U�\�(�yQ��B}>0�ӎ'�&
��Fd�C��5���)ȵ��+{Ǝ��u������ޤ0��m9����\lڑ;��Hg}ڍ� ,q�����J���劈�U���=��T���W�6u>k����#0L+)[�C
���P@��P*������/�soY�@u�����]�g#�S���US���}�ۍ��n7?J�l��p�y�n�w�� ɉ",*^3��(%���� EJP'��X��6�\9���F \6�;l����o5��[��� ���Xj�l�r�����qs�+mִ�>�@ț�Nn)e@����K�\���lgů�)Gh�����L�_PH�2���;���.J��O9l���4T��u�Lz��f���ő0����F�*��b�_�s�"���<)z�|�'�d#+�z����h�|��ȗ�a�K�D�ڰ�ڎV�f�8TW�8I���t�������F�K�r7k�犑�2��3�Y�"�_C�� 2"ot�Q\�P��<�.��:.�;��Q�x�AIr��`�3R��!���c�W�C>���<8o6��V*E7�l��8 tfmUÕ dqy.
��0�'�=,Hn� ��=��A��zI�/��.��Od����ʊ�ٝ�d��]t9��6�(-J\��i?JXK:JY�9�B�� ��B%��e�2b��HM�9\�C�WUW@­'�1έKN��x�WW�r���U����i�Fj����ty�|'����{Vʻ���ѹ\���F �����C�\�+��w�>���-�{>g_2��?��U]1Q�#�V[��]�?� �K��8� Oe�5(���&��Iy�,���2ܪ�/�ۚ��
"�bh�۰��GW�-�O-�:��#�V�qMV϶Hp>�墲��Zë[�����{]�˿
�阦�wHB��l L��7�$�c�aQ���\R%�TZI�w�	��;I�ƅrf������M�d��ͣ��A&7	�)���;$��k4���LC�� G��{�-����X��j� ��U��#2Q��n4�^�F ?�8�����Q5GW�%ESN�ן3�S@u'�`���m�^AEL��;�4����0��D$�QI2+���U"��{ɻ��i=@�&�J86	_�a�d�|=�}��j>Ø����R`��ئ'�Ę�x:*�����"t��̛H֌���� .5���-*�k��ͺ�i��AT�����Am��R��x�/�V��P�̭��L�,�\7����,z�K��<ˍ���z���a<vS���#}��>�}W,�V ���:�D�����y��z/��bws�l)�f}>���&0�H�wX,�j/d^lsIٟZ���:g�&owW*�1�mݿ�!b҃��^(����C�������'���G5ma��MFv�H�:-�B��:z��Ϛ�%}ж�Ӑ͇:����ncb!���ی	���%�m��d<0◀�ڿգ[�5���Y@��5���!�n�VC���b�s|M)'_g��~}*�� �o���~d�^#eS��������.%9k1��?7 Ji"���,�cV�ol ��� '�s3[���C���G�~"B�q��XW:��DW��͛ց"�R�����������hҞ��UXD��=h��n�>w�g~֘֍�بza�H�n���?�$���c�\m~��N�9�O]:i�{�������Q1��[Ǵ��:��,�~��k_�P�%�+ ���ȯy�De���O�dv�����x�����$���)3Q�ٔ�JO�a�l�"�og;~�>�z��To^�����7�>|cS��"r‐�T��k3q�23�j�>�#感�(T�q�k�d���j�b9Q�d�����?����"�	�zD��s�[�9&I���T�XE���l}-�w���yYu �{Bt��32��ox߉�.i�*U�~�{��sm/��� ��rֆx��a�Ⱥ��Sg?�ұ~P��ϴ�n�h��O�j�餗�;�ѤN8u��ag�L�нB�[���[Ψ�c����Q����3s���*�h+�O*{�����T'�5"�g�����U������&��G�P�/Vh�e�P0ё��/_0Ix�g���Ӥ�>n�ʸ�c)*q�3Uf�d�%!�7-�U���T�V?�:$^B<ᛈ�D��>�����/�����2��Y���H��jC��\3Eq��I�芛-��{M�1*�dG�<1ȁ"�j�I��@B#�q�(_8y�Q�y�D����R5�.eQ�d�
+p���1��Єd��Z�Ӧm�%5��y�P�
�[k�8�e�����r����p�a��\x��>#~(�� Zμ��6ҙN��ڿ�`Ҏά7�h��M�?�zg�C�7�z�kfc�G������/�ʧ�ezgLx��=�T� K(�~"�U����+��-j�[��;���T����Jge��Z�0ţ�Q�=""!}��(�s<�@ͱ� �W��U�>��w'���	���_l~�{�f����o���JVq��i�"s�;���i)k�MdՄ���Ȓ�'�v|�r��\K��ͫ�䙖>1N�.���u�<���=
'2Ed�*NJ�+������7ŵ��eU3�$�ߣ��X�TCZ�Jz�,�U6v
��@.�_0@p�md�*qiŢ�Wth}�j{&?�t�YDX�!b��	�E����y� Ě��`��Z4Kx��DU0�Hݸ��7�(tg▆�=Z����2j�/N'�Sb��h#5���q�6"���R�PA����J�A��6j�
S!�OSW7$����<b�@��!���O�$�N����.y�ߕ��ɋ�~�uL��g�		�{x��қÉ`��"$��o ��������L���/QN^ζ��46J��(Uľ��R�i����l������;`j��'0j.@�Z����6��k8v���&Q3�+
�9����^�7�e�V�2���'�Z0W�>7�ϺJbPI	̶���`��Bi��9�*�kr)�/H���+h�>=J(���1��K>���]�
Y�M{Aa�Q2�+���c�q��p{�Z͑d�ۂ�t9|�{t�=0��*gy^s!����4]K�u	ȥ4/��Tw������Ό����H�R�g[�a���X݁��,<� łSĐ�2 >#��^��6�?��p���uV���&T�$�S�dj���YG�z��vړ�^ʭ	Q9��dR��YH����I�-Q!O ��[�N$+��j�)��k�HwY���(j.?g�.Z��3+j�9L3)"0S�A9��X����qн��OJ�9�a�LK�
\�Cg]65�?�ZEN�]�.aۃA�{�>~f '�xv�y����I�;��ZU��d� �B6��9:�.����)� Q�q2�X]a-
(�q��%uT�cX����5��
Ɖ3�&���Zq�<��t䫷n�צ*kD��%�7r�[��4�	�[��㰼���J��p�⅍T!Ujk���c`(�k�`�8�k/b�O_'���i�0�K�7�E�H����qJ������ނM�*�-�bT�S�h�K<���>��¦��
k��lKmd���,�4
M���\�Xx7C����/�x�(�#]�<H�H��)lބ��0zvg���O�/-�&pQ5�o)b����%��t����T��v�[�T��۳���1t�����?R׭��n�LI����Ϟ2m���	E��J!w���ﴹQ�:,�Ɯ��F��K��[F���0����sO#c>e���+��{W���<:ϋ�����1�����Qt��l�'��^=�V�T=�Oб<��9G5� �͑�r������K!�ŵ��x��;�	ņ~~�ֻ%N��F'2}7�Z)�ŉe��G�"|����	]P,�~�{a�,	5p6VB�`c�|�7$',��� Bݺ��m��*�,N0�"~Z�B�c dY�̎P�%~��ʠI��Q���� �)�s2R�g��I>�*6bCD1�?6-A��KkTwi�2�g<���i�4�"���l�{��)�/���mz��3X�O/��A��X���]��뱘A�
��OL`r�]���0��0`?�d���o&�o_�t�gH(&�Z{
�K�c��EͩC��vȁ�!_{N���K:QW AΒq�6��0�MɞWkH	��t�⺏-Yh�8-���S�����Zȴ�N8���s|�~D�od����'$z8*k��4�*[�}��j�{�������/�f�-�6}��;�D08�O{�������_��]&���Bx���hi'���k�mK�-e��u�q	��A�Հ���up~�]i�jV�J?���[6��<.��s��7'
�躼�=r����{�H���ٷ�HC"K�%-�1��,�@*���B���/��F��0��Ъ��Z��e�G ��[�1��z�#�]x��Xf�aۦ�ੈ +�}�q%�$Z4Y*Q���(, 	h�7�,CÃ�юX�*T�s8@(Q����1��hA����D�q��|ָ#��@H�;�������#�5��D��Osa�ӱy,������u�V�k�)V���u~��$�*����y�@�D�KA
�څea5�[`1,�w���DS�+�Մ[ı�R���Y�ٺwd����Fј���ิm\��V =�]�Nc��h���v���W�g,��G$u��̱��f/P�Qu(��2����#½��s��ȍ��-�2y*�K�i�u��8F��,�B���s�P�X ����)"R0ҿr�.mv�����!�QH���A�Wȅ�9N�5�s��.`Wo�S<�T-D�"��#�.��$�����0�O��o� �Յ��ѤL)�̦���̈́�1�j;��2u���l�����0a�	�˗E�¡�{�k�Ǯ���}h�-�v�BH]�&�泬�C��<�'0�dKx$��(�8�v\rbm.�L-���ȥ��7r���	]�@
|��L7�ʰ�V/K�{�v�����_e>�K<' ��GY�]��ș�ִA����M�Z�	/݀sI�����_\C�S��讀��D��{�]�:/㜆M^��{"c��\`��Z���p�6ǈy���_�U����mfz�B�u}D�������6 �Ö�ַ�Br��]X�f���t��O]3Y����0�Ӆ[�@�O��N^�F�!��8�R/�=F���`�|�؍߀����7��@�� �2}��K$�.EN���Wm10�GzVqN̥�N=�0C;w�N�ӎ����|,���z�f<��qp�!�����>.���׸�
	�#g��	� ���v�B�|#z^������:�KM�����h�ߝ@�䑗z3�����/�z;�}�Ofu�w���0��)x���TM1{��>J�n�&)&�88n��	�u��ݏA�B
�A�����k�8�so��#�m�-k0'.uS�/��Z�V��g�h���YF�A��*^��kͅ\��n����kܳ/kPį�ֵ��:.�������\�X2v�7N���NX7�v*���7:^1�v�YB������r�49��Ih���"�2ŭ�I�:u�� ]��c��/|@r��9#�ʄ������&ΕX`=�jc�1ґ�A�=�?�/7�
lO�0���0�ɍ�֒�%����ޕ~��&��P[�@c� �A�� k,��]|�x4uq%�}=Q�;֍��
�#�,Yb�p���b�cR��?�������z�
�C�$1	�K�q��$��R0�l��V�����\��#dC����%gSw��il8ޟp���q���w�sշ^T���$($�k���5�30���)�9�,��Cv�`4�8]���0�(W�>����o�l��n&��N��t� /��$\�����y�C,�R���,	��+�jg5�ޝ�|����׈>d��nR�o��J�jkE�nXesv�x�_��C�!��Xr
_Ѥ�%�L��γ7��(1䭼�K�\5�����7��Ա��Me	0�rCz��mAߐϛѥņ��������D�p�& <=����7l�f��G2��zuQ-�տJ: ��d�>������í�A ��/1��Uh���3wi��w�)�o #19�ߨ�A{��'���U���M����Vв�4���������q��Ƽ�BB��E�5�@U��}��6%
T��W\����ͱI��W[��A�	�=��e���f� �Z|]��1{����{���m)�aǡ4�xj��R7|�u��	3�j{��;������Q��/�%��� �'�ꩬ�{�}_�����/q c����.ɹ�����i���ǘ|ڤ>�l2�ji�E�'�x���Ѡ��N\l�����u��v��!�02׺�$V�v��9������f�V%�GubR>`�y0��k#�3�D��չ������U]Ag �1"��"[~��y�.�ύ����K6�K��/E6�V_�#�x\��p��L����82��Ն+��p�w�V3�Vj�8ګJU9���d0��.�Ė�L���Y1��l�3&���[������V��	��`PjU b��Whrb��2r��F�wt%�WG����pü��i3k^�4ќ���USܯ9G�S���M��W�Bʋ�Է���z�/����(�,,3g�	E]��4�Н�L�k�@?��!�@l��E)� l�JMJ�b��}�5�kO�@�#�B�^��׻���/�~�>��/,�cvQ���<�.��*��m���`Z�"�����*؏�X���,E� K?^n�h)�����f�o#��1�������^�qմ�ҥ-�{�S��%�WǾI��Q���-�ִ�ٯ�A,����D4���:WnX�W;<����+��)+��x�w�j�s;e���5��|6</K �~���3�r�Z0��PA#C��R�� ���`p}����pE����<��V����uW��ПI9�oZ;j�/<�E�EJ*��{(>h��V�2��&�}�6���������S�ٷ��$���S����[�r�����U���;	� �(`�Y҃���*�^�By���(Ml���V�RW,6r���ދ�T�c�>�m�V�{pB���@�6���zW���KľD��9w�M)���>��@p=��\s@��?�~j�0�:IC'��VU,�q���9r����yIN��7H)��ZEbw7��
�l�Qt��E�v|����Xj�Ô�� �Y��5Z�tjߑ���/�S$�v�}js��ūi-p�&��� 1����n*�Ё�NI1{�Yb��)�Z����(�p���^��G�}�v�:(l:r�VY"o�����j�T��������Ɓ��7�\.7�I���a�<���1{%s�43�F
�*���у��Yc�6hŎT�Q����F�ުΦ�f��$��{"���> �[J�?e�J��M&��J�7Q	�=A���,�*�wk�R������υ|>���E�"���I��v�������$�BC�.�|�=&Y<�D0q�P��]����0��6¦1��?PN�E�8�q��S S6bp�r�T;�L��2�z(I�T�>��,�؆�W�����s�¨�,-�Q���s��j�.27���K�=�nLQ����h�i�r��5��$�ړI�{�T�O9�%l�]!�*�+5ӇH�e);�)!$�n~`����_$S^�f3\0�$��eyN��z�ΛW�v�OǄV��z�e���e�x�O����y%�k���5{Y�q6����/4eR4Q:��\&J�,]��s��
6F4��Mb��[���봽�cF��pk ��~,v^��Z/��	1 _ùi��w�DY-a��9p{�aD�=V��g�+<��^�Y�JzOM4���w)D��<9�Ǻ�E�	�1�J!�s�D�L)��/�ਟ����%J0���R���q}�u������$��G= _�95�W�m�E��: #֘�+��Ȩ�%��֙1��Yc�"w�4�v6���Ch��XZ)��Y�9�V�w���� �ڑK}�ݡ�gls�������a2��M#�Yˊ���T�K��o���^X��q���r���G^�a��]#��XyƓ~i�BB��1\�89����Ӻ���j!�:Ņ��N#J4�p�&*��-ƽj0���Fq�ｧ��փ��)B�w�Ͷ��))XA��)�&)B�Rn�Rm�~Ӗ]�a�}�I�#��7�8�뮢�9*W�=Z_����X-)��omw��7Z����/A��o�v�B�o�R�&R���+�>�a0���c:~bq�(i���=Gٚ}c���er��y25H� ~�]��T�U�4�ğ�'��dݙf��n�	�O�(��S�P����+DTS��<{u�o����I�ZmK㠛��_8,B��$�]��e֗n����Ym-����[��cJ�%�c{�jv�F_1�cc�iM}���6v����W�LjXN�O>��;���i����K�x�N�Vo9�9��<�a~� ���yHФ�w���փ��L4�fJL�Sl�/�lh��(9��k)�v%�h�,��ٿ8�+gnL6��	H)�6A�94��p� ��]$�S�}���7Pw��p�o ��p��5{L��sT+�r;�a��9L�n	�47�?3�J;C⣚H��I �f� ��=�q��$�]�ZZmN���g�ͼ5K0){��xK�_B�H]0.eyٷ��V�ۮ%��N(D�|YU�ѩ�0��ѷ��Xmy�GP���I�[yB5�=�Q�m�������'���`$�'�]�X�H�rN�HF0�����)e,s�'Kk(y�3]GP�|T�í�zL�9��t�?SW�;	������6M�~��#Y�B�U@a��c�v��<!Ȁ����q"0/X���p���>(NGyߌ����~��V1��q��|��y"�b�Z����6�� ��2K#�_H�\�af�-�슮�\5�Kڂ�7_�u�f�"ѱ�#7��=ƴ!���:���
�ܮ:� �4KN#�)��x��qVd��VnI�V_�{nX����^ԟ�\����2@'5wI�٤*�Wnt-��!(�����KV�!�k�XG����C��dX�-��2'�/sÃ�s'18�<��it�d����}��k�9��[���}I¿���{|�!�1�瑍o	�:#cS6[B]u�jƀ���:"g�*�9ap�	y��(Ǆ�$�E4�G2�IE����H� �fY��(R�XnexN�,�$�H��"G���U���	@���ۃ�@g����zʹ��z�G�-0	�d�}}�e�J�_�|�"(V��~�/o��¢N�&7� �J�ت�C��o�C˨-��s�s�G�sΖ��8�R0;%��#f�����=i�扚P凓���g����+���5O7�ނ����%�|bB�*�
�/&1.�l��=�A���A2���1n37%��te�B��#���8o	�DP���/�����ױA-�l�����uo0���:��Hc�7�����F�����C�
�Yo���f��T^��� ���r4�awA�UJ3@��'���sl6uA���61�dq%��h��T�癰.T<�E��%�]��O�c+���(H}#�x_
�fM�ӥl|
���,�\�Z+z��7�?8��H\'���s����H�Y�0��M%@�.�Wh���B��w*�کf�L��X�f���QfM�Ǥ-��z"�QR��o��8��u��{� �e3>�Y��i
#,�KG�0
ly(��&Ce�'���������"(@n�Z��)Z���أR�55y���C�ظ����ͺ�t����ZC/���������n�M�Rw�Z)!�L�Jһ�:��q���W����+���.�e�ӣa\�h_CQ��.!e��
 Oeu4/Ь�|ۼ��4'66�16e�~M���6QF��Ǫ�\��Ȓƀ��z�?#����0���$�P�a�@��%K�q�eҐ2D�,���a�o]]_��g�����+�	-i�=�I	��F���-OXC=�gn��x0j	B��O76��c�6�"��=.e3��ik�]����J���?�nza���7�1���ח���/o:X�'C�i���(	�_�.�U�2*ɹ*CF�*�	�C�o�MZ���;z`8�f�\�a�
S�G(j�]�F2��9��O��#��7�Fq�WH������h!7��c5�g"�ZN������oo�&�k�:�$<!�MR_��L�D�x��vj�vOY����L��풹�u��@;'c,�q�JhI$U_���Lʐ������v��̿���=no�/�6�Zs�Kn#g��{��,\#[����v��=7k�X�� �{���ޙ���&��� �U9 /��q�0��8(J�t���*԰`�E���6����~kU�҂�e=EW����OL��!��I�1�{���q�L<��[���UX�u�u�S'�	I#�*��O|5����Y;�V��+&���HI�\{aIפ�6ՠ����`U�TF��a����mAG�ԃ\K)�G#ð� ����g�_`�wɮ����S#���k޷��9��T�(�=G�"��an%�y��ΔIf'���g��f,�tVX��{3Շ�P��;���8�u�{��h@�cك�i�8#,<[΢9\�E˘�ޙ!��8M�z��%��D� �jVKq��n�0΄��H1�MO�����:ئB�l�m�y�U�)�B�v�wf����?�F���9:�B�#�&e-�m��L��~._�A04;Y�#�n�;���f6f�v��n��5���z�Q��RO0��gN�����-����3�O�ѫ������e�󄓹ئ�F��![��E{���/RH~��+k��[�������|�lЊ��������2iM?itP�I��� ���$Aͽ7��ڛ3����,̀�"6?����&��Jr�I�BvL��1S���#Ϛ�;ۚ4;֎��+%RY=λ�J���%pI��aċ,^��p"7�����lfޛ]���؏�S�SkK�:�d�Εjw�X�W�F�E�ƨj��*��&ˤ�O0N1A�F׋8���*�B.�a%�DT�Ckg)ڻ3 ��:4
�b�Ax�#�wق�		� C�ڑ��3�����x6#�8��l��+��t.n��e(K
��K�	���W�#&��k�MJMq��ǳΛ�a�;gKg���[C���y�5pR�G��Z��WGx���]�ސ��
����ɜ� ^?��ĶY�L���r�:5
s�'r�G��#�Dzz0�W]O(���V���Iێ�߿I���f�K>�=jC���o�A��mcg�����#m��}gW�@tF�5b$8���˼���[Ȥe�|NR2�	�������p�}E����gR���a�W���u{�f�^f��(H�s=��
�|�!�c��@a�pb��M�0:�BQ&x2)/��̈���	v��ً�w�B9th9A���b����5�Ta�h��k�� Ek���QNI�,&fP=�'{f�$eu4��a�`�UywU"j�-0�މI���= #�`�V��s�����bW�ݳ��}O���K��<'N��R�#H���Ƽ�'��^l��u+d��b��1޶���D4S҆�Y��yaQ2c���r�5���A	.W^��Q���{���QL�b��L�rR���.�~	t���+y�撔��'S��#nvC��RS��E�C[Jxl�*+"!օz65�GtRBi$r.:e��;��[WB�8~fG�G* +�#ꖕO�W�P�-��ro�-���x�뵅��+KET������r5d_�Xv�x	EH����-W�h�j\B�yp���}�)�Mq���o�uu
$	�FLD�\�� �ccV��%g�A�ȯ!P���B�y�~��LW|s/Se������k��؋�sC���c3���-h����������z)՘|�� �謪eu�pl	O;�Ly���a��U����Pv�񺀝�����c�5��r'҅���� ô�������Q��0<��I�Le�N��@��j��madNL��(�~49�8w}I��c�����0r/P �@�ə�[?F��XJ�⺛(3��sA�-$x��0���4�5=�A�����ΠB����>Nڣ���w�U������Ct��!������8���4J8��@�\6�[Q&Uz

w�|�Ϊ�)�dkt���V�z[����9��s{��&ܝ��LX�mH��]#�+w�i_�r�mB: �o���e�w����?��+��eNI6
��	�*�Dh܀n�B����XX�����Xy�V���t�@ �m�Xt���@��ڰ�}d�u�^~���{�O���q�5����1���~$id
�;��L�c���d9 �b~��9._2[��YB�W�V�x��ug�h�5K��L�o�7�ɳ�#�:61h:D	�T�2��	BeW��U��#�^B��"�B���O��}f�M��ט�fU�*���w�I.�H�v��}m���k�Zq�m䪯���yR�RiDb�n9c�R�M|�v��U�+�D{�*���5M�S
��X�ħ����S����H������H� 
����OW��8z|�$,$�Ъ&��ʫc��%q|�Sy�+$�!2�nN��̸��wSa�Ji�RKa�Z��h�ɨ?��`��s4�5x+@9�Ǩ6�gAI53�i덜��Ez�)�WK<�������r|+<�Y(�&�.
8��N#5�䊫���y�rP�mo�{d�%��4�߲w�U���)��9k50U{'lK�!6%2s٩����;,��>����XV��S�*��ҟD�D�R��f'��S!A�L��y���kM� ��	���h�a�o��O�t�k���-�oMod
����+��
a���(��Of�p&rP(�+�{�m���F�G�tq�D�+[�A>��jrN۝i6S���x$���n��?�7=�`W�;�ĞБ'ρ��i3-@⣬�o���=:.j5sq6?6�������l���[�ơ����k�:��u�qc�-�A��- �O�/Y��E�����xI�H �ܖ�>AR�x���^�5A�xO;t����'?h��^	&��{���i�BR{
��D�^�X�
�Yj&Q B��4�b^�^C	`�~��q��¶���f]�OD(��:�R��6�r��K!����X�8/�����4Zϰͱ�\���k RH�>��'�F�+C��2"����j���? ug�w�m�{,:�>��,᙭����h�!���Y��M���0����I⃆�xo����\wkمP�)(� .�KSp�n���k~��ti�/���+*�����/��A�7�`l�CF����5� v�+C�-�e�\#����#�􂔀^cFy�J�-����Yd�O���e�t������6��U.@�n\���?�<�	�b��16��'�,�$H�M؞e=T���$x7�3��$�h3r�e�LK��X�0��J�=�N��?DT�,��f�չ1�$��U�!��!��pg>��_5=�2�I�9h!6�;��Do&����/�>��@���h�`#�/���L&6#�e�6T�B$ZŬ<4��P0JT�
�[��VD�웫�<�ɫ(��[�,s�ޣ'���8gs�];AwA�ay���&;5��;�$���p��J��M�\��t� ����55���ە0���HV�G=��!��(�*�ҽ,
�
�Jq���"�Q��z�TN }N�N���3�ܙu���Q��4ڶ�&J�z��W���\��-h^����#��x�&�����<#}��0��,�۰~������SES�t�>@�� ��?u��W��-mw	U��˨d�Y��؀ҟ�L�O�[\d�W��n���(T"��f��/�5���׷�EEA57<��0=��Z�Nj�Y�� bn�7B��D��#�_����5M�>Q�ʇ�LP�Ȟ��G�� �Wϼx{��v�0E	�s����ІL�'(ۑ�X���W=���T.�[XW|�6/V�[zZ�0b�/����}��久����6me�̑��e͈Y� $��K˻gM[38m<>v��C�v�c�P�8�>��2S���"�Lz.#�Q�VX�m����V^_���$ۯ`4(�<��U5�>B�m���u�l�VD��X�uZ���:�y�,�m�Y��p���\�����{�����m�[Ey�K�g�I��;�1�� �tr��*E(�2��^d��DHH�R�����T�/�/3Y�62$�Y�B�X˥��9�P^���)�:cZ��!yȯ�c��Z��=�=�og Dh-��1_�tj�����3���SWR�x(�4�)�6\�:uh��R�(U�/�@��Ì�E��T�t��L �{�7v1�'�Ю�:�	�#���v�S���<F����b�����p��8r���d:�w��
�w��2����7C�OĦ6�Ɩ����	��Y?�-A�)M9jS��k�ZV�O��qs��ZQ�"T]��X�*��tӴ>CR|vOΦ���^�{�A:U'bG��w�;�@�Wð/y#fl1��	��?����+>^���Μu��	�y}/����������;
#�xi!悃����]�=V���jkD=�X�
���*$���&�^�"����QS�����N'6�K����+��A9�Yp�Ϋ���H�WT|���WZQrU�3	\ Y-1Q��,`��aS=�p����ٿ%�X䕞f"cU}1��g(�	��T{�]j�\Qޞ��!rY��S�2�3)W{Ԡ����|?:�yA������Te"�X�(�A�������qH�HxxI/#se��f� u!7��^p�0��~�Hq�[�����FB��̌)e�l�����-��:�a�|6<󁄻�:mTA�U��,z�Ya/�eO��������%���I!=Hs*����Ȃ'��v�Z2p�V��1>�O���b�gI�3�]{�,%�@���t�Y�]��)e�ʪ"$��,}���+��=Y����[��ث
71������.�AC���� �#N�V*�Py��
{>%��#�	���@��D�:�i�p�8�mx7�m^�6��/�LB�A�b#�(�	���0O����,{��H�q�M�Yl*�>Lh�n�����1�+��i�M?F���Cl�����G��g[u�(�5S�|��Twx�؞%�8��q����rp6���&U�z;�]�Ð8��Vp��o�/�J���v��l�3�:�M�$�t;��J;�u�����Iz(�������ۣʞ�x�'���I��9�-3H@z�՜d`{g���ce���J%�bQ4�ND*��u��G��w�En�s��'��s�(6�N���^��"9>��]�կ������ɿ�7�o������{ג�e��_@�@����]%��� ��*��H�!Ҟ��
��A`����]��C5?����l�)��6q�!
���c��--��e�	������I�z��+����>�듗�#�uC�&�+΂� �f�꓈X"bj����;&�E($��C�����s���K�*�ut������(pp����B��;%��qK�M����;~;4���daI��[�XX8����S@zT]g�;�@'kar��Z�c���'�F�0� �;�,}Q��77^���W���D.�h��bq�&�*L40oKd� g�ߖ�D���	<r�p��
��L9�)�{�����9�q%ס����+����f�<��r�gH9�>I�7׉��i:���`��H���o2�N,|�w�!C�c1�s�Vixq_js��Rb�!�zyE�k-Y���i�%!G΀����0�Ht��D�vBaa�Ų�ٱr�Y�S
WP-�8�:�������D��χ4��'&�-�kX)i�`�=�����RZ,\ʗdߦ%R���<05ؓ�A�EdJ��k������F'�^����tR�w�^��v���\ ���)�d��(T��˾o�L��[�ʿ��_m��|�q-�H��NU�#�=l\jOL���]#�OT��j�@�"�5r($�����S%ˣr�=�S��CY�=���G��+�r��%@�>-��N����m����it��XA��5w��"���J'Mg��WɈ��h���D[�ۄ��3��������E�Qs�7巪9��JЍ%�{��c_�>Hm��s�ˡ��Z04��$�: ���f��6��:m��'�e�	�o:�\��ʸ?��~���F�L�֍7*F����|U���qL�����͢��7�9}<MQU5N��s�]��<���U��z��h�p3e��i8�Xpb�<�)��W�S�R����'@T<w�v�R��j�FH���u��JY���ĝO;7ÿ�?Qhb�f�l�~�)"��'=��D}��js@�A���~�����A#�#�^��d���ִIiO��Zb�l��x�5��y�洴P�����������n���1�9!�ٓݣ��]8ٿ�튒o��yK��q��i��1B�}�!�r�4VixNeМ�s2�9���4����-T�{��g�5��;����x�]�;�k�z`Y��06;�Y������,�c�:����O�1�5�jt&:���m�N���$2�W�}��s��Э�v#��sxYo�����J5�����Œ˴>Ϸ�,r�^C��9�ߊ?�bK4��c,��L�h�����ҼNs:N�~�0_�Vްœ���њ�׮�ꚯp�1��z6աc{oX�j��2BX�p�M�!0�U`�4'���"�t;l��ɦ��'���H�	�q��a<Dx�����z՘���ɏ)�������`%P�!S�t����y��@�,z�:N��U��Tҝ����=��c2"?r������d��[O��р.F�!��M&A�}d�s��*��N���l�Q��Aw�E�[�e푂����dާ�5��N�ȑ�������9̃��M��� j4�?�2��(ex�M�34��#x4o�l�'I���Hg��7Ա�b���͐B���>HS�/��
ݷ�a\1����E�s��91)ET�]:6�ք��b�}�l���s�3=
��-�����s<m�̷<`�|:�ځ���h���?��������,��R��HjM��|�B��G(���˦ PBC���E����lu��u�[���8}�胇����5�
��#����v�� Y� v㟒&v�?��B�nѽ2!6�D9��u��=cd<�����p��6jIg�x+��5T��#{���!晪�9j�;p����&,�(�7|P���澨��l�R�޹��ܟ��xћiF�$�c��+�Ã"O	��mS�3e�&��ip�D�%��k���x�;���oR�CJ���!�֑���|���W\姵K��r{jd��#	�����}kLqMIe!j�1��A��(�j�[9	��>�}P��2y��ۜN��)B��a u;
j���x����_�����-���������$I�����!� ����-�.�B�p䑖�|�=lh�"{�KP)�tz�]L2͂K�	K�[!���T�{.z["KDjXlSr�[�t>6��ފ�3���'�&<�0Y���->�?u�$�|�\z@�B?�O�ӻ�5�şR���\�Tς� �o��:�����_K�D���� }��H�W!KC�[�j��̊͘���k?$�j~�HT�<,�i0T��/K���W|�FJ�aW�hHyVZTʯ��<[&�9��I�w?�"Os��h���������e�٨^��L)a]�}�KS�)Q�bO�yD.Ebݐj��M���?C�՟,���!z��^=G�����N��?9&?�%���4��~�V�E�`��D�(�Y�C�m�Y`e�YU&��"���#�x� x/6|i���FX_�͌�#-� O���Uշ��L��R\.n�-�H%&f|��3'����5i}����'|��_��i�S�\J�)52Q�]Aey��إ�K?���J�>�^�+�9+�}5���H*�
LQ��� h7�77���j�F�4)_)�E�S���ע�6�6���B&�>�M.u'�TR
�*;l��ӫ�*���PD��H�@�C�,N~׌}�mH�\�>�+�U��8�[e�l�Ѷ�:&o�d���A�B[�x@�ݑ<�(���y�C:ۓ[q���\��ǘ�Ѩ54Cՠ��@+_x��}y��VN�K߆�����h���afK���\�&�GC|@��j��`��&Ř�m���*�P��;��ĺ���U%�u�����i��T����fS�w.=����$L��`��G@���\�䶘��;Q��Ȃ�kp�S�¾���;�;U�.D���\�,����;	����Nƕ�7+r�i���6Vk^��2�CIKY�����+|^t�o��܊�x� 	�ķJd�]�j�҆~��dS�@ �vWjY:�%"���m�� _�Zl��=5K��(�$�e��XW 70�_s����j�J���)���`[��U��º�F��CH�B��qh�����\��}V�$��2��ˣ1g�z��]����æ?,�c��ܴ4o����0��O�-yf�𨎒N�∥U|ëu��������Q�#D[� �'�����&���=�4������Vf��}� J�O.ދr��.�̎�e�;>CR���8�YYؓ�Eo�t�޸.;�L��Ѿ��:n�v.�z���.#g�Yh'K�x��z�Hˋ�B��"�2�'$�>�6�����>�"�� F�p��� 吙���.i�����֠zTʷ6缐˵�)@�t,�!��`��Y�pT�8�K%*�,�Ƣ�ѼW/���P����X�8<FaV�؇ ��,����ct����8��e�|�$

�!�<N+���u����8tq�ұ�fVM&��2"��h1c�����boO}>~ۣ�α��&v]��(�ש��M�wOF/�Q�R�z�@(��`*e�	7���c��t�fL�*��#9�͛��zg���Q���o_ӗN����O�EW۸�=j1�:�g��sƹ"J�Q�'v�ƒ}�X.N���Z��J�Q�>����D�.�V�3��K�T	���OZz�O��y|y�Gȡf'���4�Qq��@G��h�<���-x�%�z�B�'9B�]w�!T��x�����;*��_�H���3�fMn�C�uAr6� �:��_
�[�p㘽�Z����Ǎ�u����5o`&�n�g|���@��I*�%Q��Gh+��֍�D��F8�N ��^I%�X��?<��.�vWm��b�6J�f�إ�P�۸*u�s��-�%^-����H� �ۻ�@��O��_e��7݈=��~�!�gR���>�HJc��F!Lz���V��T� �G��(y_��MZ
�ס>��8��e&�#�}䕟9�-B���]y_b딾�����1.ň,(��21��Y��H*p}񏽿�>!���F��qUmY��q�)���/�$��d5o�����s����qQ� �e7�ؙ�aD* `f��r#�U�vܘ�ϔ�<���;�R�?�Q
F`��T�5A���φ�Jcp��<��<�98ѠR�S��8Ѵl'�7=��\����Ȏ(6�X<����Ð�ǈh�^���{y�����Ԅ?n���%���)�r�� /�d���Y�`��c�* Sg��%V��_l�3�!6� ?F��)RMi�W�F��w�[m+��Wp삊92����� �=�濛�ڣӼڙ��t�Q���2����Y�t��]��~��d{G�� $��yvE��˻�����t��+u�-�a� }���_��cq�4�ŋ���|7����M~��� ���B�g�R�ue�> �9��3g������v:]m��&�(e�}���@�_xxW�2�#sqVY5��&Ogޖ=C����a�A�ߦ�"lC���K��J���?����>q������x��;K�6�eoa�ڜ�c�5�-%e5ݹ^���6]��j�t?F��ֺ݀�^e��.2R�I�\�7L!J~��*����y?)�y��B�Q@�	����0Cxx�oa?��)]sl|STI\�}�	��PY4(t:�~z"s�/�c� �ޚb@t�ڲ���Y���d3 ��ɩ[˹���|?98R'�H���.��~�����v��:yc�`K�a�Z����K���ȏ�1�-+�K-��������ݧVÇm���÷�_s���\�U���4hk/\7�l���1�����zёfO`�3���"��F�Vv�u��N�lR���1��Y�U鼪TwN��0�H�i��{��_���Q���i��9�R}|��Z��̯���h�sW���[F��3V��<Fg#�~���A���t�K8Q�z�ק�r0-����\���s'�@�nKc�a<�?�_Ȁ)��?���lL��R�N�2*��.̼O�[�Ҿ��pHݮB�l�@ҭ9m�Mʻ%N�4��|4I����𡘼3+�4#�O�TsH��^/�S���.G;�}
+Y�n�ȥXF�{);�Lm2���5��<�R�M��m�x�v���S!
�XQfl��(�2-Fv4,j�c�M�cǖA���X�9���4@ ��ERG��46
1��f�>�v�0=-5����A�tX�"هu�֍f#�E���R���/{�����?߷��>�BCq��/`7:�D�Ȅ^a&�n;�o��mCp��v�}^�+a��;��v�PA?�%��Y�M���协Žs_���l�q�d�f(][uYs�M,��t`��0��T��K����nڟA?��y�ó�	�ax����Ȉ�IO�B�ЃtX���W28z?]���5��[Ti�] 鼟bl�8ܷf�7�����Ӎ�jz��m�t)�����5b�M�,G�-���We��#��b	>r���	�^���ƜFG��͜V��F�����e*�i�}ou�M*�|c���Հ��+�"(P����C,�9:�'8N�A�<�W���塟�N�vO�O�����2{�QG�]N$������N����bii�IFZ*
���]�xZ�D�=lf����XR�Os�2�Jp��Ƴ��g�i���/˜�&�ӑ�ǣ�q'H]�2��~�J��S�6���vy���ū��g���\(�G��Y����j՗tz�\�2��m�rgzQ��zy���б\�����2�˘6$�H1��J}�����7�ϝ��͝f`�2������"�o+���m�]�����C����L��Y�I=ķ+���_��u��%a�cⰳ�1K,K0��c(��֕xV���;_R�I��gX�'����n-a�z�@d���rD�7�	U�mM~2�P�0T�|��E�%�]���
�.,_Z��I�b�����`P��&E�}?e��3�#�IT?��t��B`O�k�`��J��'��՞%���O����;x1�<u��rC\�DaK�ր��5]HԽ
����J5�h�t� X�;�|��/\�s�=4��ٖ��6�+/�aO���ڤ��J�%���-w��I[ƾw�+LG [B��~.CX�N���A���8�!��u���N�0UM�zzh�E#
�����V6s�a��1.�����,���\\�^r[ül�骥8s�֏��$\�\ �	�e��Ƀ�|H{�r��F�˒��p���+�r��]�8J���Y�E�����R��*S�ץ��}`%qu��1��4o�,��f���pP�
<����

�at̃�<�{�N&����^�!���/;4�`P���4�&ڎ<�.�n��I��-�MK�0�?f�����~�jޯ3h��#ωZ��[��H�D��>���g��a ��m1�-؀^^v�t�2W\���sY��R���s���aTLĳ��T�Oo�Ae��b�?=xv����@0$��,�C��ffu��Vaf �ݖ�p<�%������{ő�E~.R�1B�N�v?�W���[���vx�iW�E��bB�[���k�A�&�4(�c�\��`*O�a%��Q�L��IC����+��������(P�CS�o�Oؖ=!�rֆ��T�Co�:�ڀheR�W��p�^4�L�
�s��.ǯi5�^.��L>���F�/$Y��)��Fl�r�Y��uG2�˚�̨��]�@S
Ӆ���;��P{���7u �]�D�i�8#5�5�C����z�H��m��U2=���.��������L�
�p(ڜPf-F�Ǜ	+ 9X��W+~_M�W�r��Y�x^nU]�72OӼ!�'%��O��	sXd�E�2����L�9���M��ʱ��#��E�P��u�$;/�/�#Z ��o�cg8
�E
�<���PݣA�MT��M��}�d[ƛ_p ��Ή.��HDMWs�%ɺ���[�_��u׈C#"�3��bZ�'R8~��$���W�U��F�RA�a�<$�n��z0:R���hwO��0�� 1I�t�/�G %j�Ű� �qH���}���a�#g��)�_l?�;Y���=f�)��S�U���&+�5�����w����(������#�+��Qq
ʝ���i�#��w���FS�t�Qg�ӵO��=�K���\���)Z�]��ϖ�5��a����-V��3���!��L����!���f�ݕ6-��b��>?jze�|�J�}�裱�d���,�@T��)T��ʀ��Wά�Ai�%����FAw�I��!K��~��G����m�3�ڀo y.��d8�Ε5��U[XXC��x���
9|OnGխ�J�:P+�닭���k�3 �f�Bl�ƶWd�Q�D�9���?LV:y�a#u}*���~[d��y�Q�4�O��oG%���Y-!Zʃ�#�����Il�OU�G�G��z�;T���L��,�v��?uY#|.�r��YX.-6�G�5@a+D�ѷ�p�f����b��B��ѩ.�%���Yw"�Oק���BpQ�.F���$6"��bVQ5y4��>���J�G/��%J��1�\ڡ6���]Õ��P�M�ߧ���}5��?����u�^F���(����k	F�?z��ڪW�sS���`=�E���F[B8\>c��.j�^JB�N}M��x�,�3W�7hѪW�KY�����m��&ҍ�o �ms�Դ���8,�J�!�-��/���Ծ*���ƨ}� ��!ylx0|oa�R�cM���$�r�,`�l�$�c^f;�;�]F�dF;�t�����;)�o{����zx-{oj�/�YS�0:>��MH�e�(&)��$3Ӻ`˯�N��C������>��	�%'�Z'a�mu�!$$V�A�Q�p���U1A���^8�S8����Kzn���4Ky���zB	���=�Rd�]e����E�E �h��92���O.d�<�F�j��_�;~��(?T�ي��]�X� ���ǭ���E]v�*�m.�	
�t�����p�_�x6�=X\��(��j=�xJ�ɡ�$fjf}�~���
ҿ�)Fx�/�흁�`inُʓ��	� ���r4���j&�	����S�r
?��k���b}���:K ��9iD"�q�yCi�#��jI�
b{��h�f`�g�<�rfon�6�,[�Y[��V���o���@܌�fG���M��E�}J\��c�W��l��煉}�՜S��%�q�$�Y1I�a.)&N���b���������Fska�+�r�H�7�:J������)n���>D�<{]#�e�Q:]-�[Q�c�+�wc8�@�=���0�5ݽCA�j5w*�d�����ΐ�������xHY�=�iũLF�CwX��V�#_����}����������!2䔁�|>t)�h"��+�q�G��sj�[��'yR��������kvO�=/�f$5��X=�������&�ۛs&ÌJѤWb����abU.A�
Q�[5���L��y����8W�O��P~W�n��0�`*؍M�`��w0b0j���7�cD(�!�ե�0����*�JS�҈�s&%v;X,l�@X>��q���)���Dsb>l�ᰗ.&��ꂬ7H�6)��쩚�ڈŠ���	O�Ř���6+��逯��IG~������J4c?nQ�����VU��b?�X� �̼��@g�x�D�DT��u˂҄��I�,�t�e;Jv���Z�6�8jEш�ռ~&OoʧrS���'�.�Z��7@�`��W���@E;�<x��Iw�Ԣ��a��6x�j�u$i:O���{�Mz�D�x��V汨�cB�l�>�� ����P��mU�y����1MU���u2n����; ��,#�K�����"��/ ���	�Y�;�T2���+��C���qR�a��?��<_������C�[���ӳ*Q�k���Ap�퀵�U�e�i9��$���-W�mD�q�f����%j�˶p��N���ĭ�L�j�S�MshR�M�Y���C�x�����8�/��-��_J�=w�o�c,]�J��O�Bk*��)�%��d��K�82�X5'ǳ<��?&��`���k��ѯ�U�f�F]u���}[���%@�C�~.!B������	z�����
ډ�����'�1��ח���7cJO�)ɸ.L��@b=*O��4�;qY�#RS�t4�nNR�_G)�	e�L&1��F�=�:������I~aQF�����}%���TM+�x���}�{\a[�S�t�
����<g�2���H�c� JIqԷ;��'MH�Pn�i�(��Ș��{~~�KV���x�nF
2z)�I�?�/��(���B����n!��p�OKy���"�
��M�uW�6��Ug*��x
��ΗQp;�@r�������;�D� �	�#%��eI�'Φ`c�~`ә�lS��.��=S�5tJA܁^"���6����g<��0�	�L,*�6��6�W3����5����MƝ|A�2aB���ٷx��t��4�X��p%�!^����8����
��;�	��H6e�7�ر��iZ,!e��-p��!I>r��<R~!!:�i��J<k�����!�䮋Ws�9<x�lD�݇	;�޹�Z	?�6�������~�\��
Ɩ���9-��F&�A��U�ɧ���]쉴��v��77瘩H�;#��ܖ��$E~4���9/���b�Q����S���Lء�4�5���.5�s�xQG�N` ODM�@2+�Xu�R��fֆ6���>֘N�t�����T/U�2��&"L�l�ӷ�%+ET�R�l&Q/�}���ʔ�,\����;��H�Z�[s��+�����6��Vj�E1��7��]ӝy]*�.�.y�{���h������E��ꖆ�Y�����)A�*��&�ﴐ\��8��??�U݂��{{���?Ώ�BQ�gX8�$�P��<�O-\����?�H���l�h��73UL���w�5��N9�I����]5r���#P��$.��*��BG�Ú�NZ�(��B�6�a� ��yX�8\�}�x��Zd]������d�K�7p�B��r���"�/~_�'4+���C#ϓo�p
��(���ݠ�Yrn���i���vc���EWD9�4�(�}��L��eJ���~�<���
�/���g�@=^��@1�4�T�l�0z�z
RgB��?ؙ{-���f;Jĵ*�=P�g���mz�#�O"{b+�L�<�Ճ�c�+`-F�0ɍ�i*5�9hden����H���,Gh\��X�������Q�a�?9P$b�&�,��nq�Zw˄4�rBm]zۧ����u���m�$�M�7\w�;㴈dU�y���%z�5[ڈ�'��^�,qs=nr��%��AȹN5��j(���qѪ�����WK�Ecj�(�Rr�s�����/E��8{&B]�����i���ʕ�e���}�y��'#�\
�kĩ��ؑK[jҢ�n!���VAY���'�l�i�#-���&u�C ��M}g��SW��dD����TvBP`ۀ.�]3��18UO��
������*�#���%x�9ő����2�[���`�NW�%�Xߢ�ɟ"�8���+E�4B�!���f���g�<v%g�w�k��Z{@��4dh`DH͟ �#�ͮP��|pqPY���Es���J�w�=�~�p~*�uB~M�p%�j�K�^�v{�Y��R_1]*6]�h���!a��tP-��G��el�?w��(�N�/��]�e#`�f��lT��\���|C�(*��@�,xm�9Ww�`�8hz8�d(�u%�[M
?Ef��>�<��6I��8�pH��n��vh�9X�� ���<��=r��Ѡ�a�Iҥ�T0tI�7���'qJc�Qޅ��"K���������"��v�#�w�F���6�����R5vU��pM��cB�X����~���<q�I�U.{U�3���4����?1�50y\��(�-����ZȆs6,]gi#����?_>
v�bsisp�J����S��� �[Cj��5M�[#��
-1�U~����y��� :�2�����H̴U��u��~ثg���|�f��k��z�[@�ՂuM����]�o_P�ȴ�d-F
�^۩�Ye3? ~�4�f�&$j]����ۏ|#Cx��c&��4�hU̘�,�� [�m48�{�n.��n5��%KO�囬��uSވ�!~{���k�ǔ����*X�����u4�WQ6:v��vG�e-)t��C���i���'���E��=�kI�a�2��R����-L�}����V?���~��i��u��L����h5ht���!+)A��*l٫Q��������ۓ�뺸y/^����>�7hK1'n���g���|��7�24���v���Q�ra<&��$uN��!���'��tdr�h��@��|�ϻ���Z���W���ɛ��>������l��g���Kۇs�d&��[#����P��I��I�I�<���x�%�yR�]�_G�K���xcMԄ��L��NG�Ë�$�00�H�C��Ծ�&G�r�P��Ր¥��֭PK��X�3zYV�%ƑZ4������Y�Ҽ(���8ZcK�+������r2
x�����n���kmtӣ�V�24�B]�nJw^2QĄ���!��>f����.\0�>6^�Sά@Vl�F���*w�W�j�D����"�aո�oHk��:�Q`�rK�G/��}1
��
��
8�>:�̀.�:K%�O��E\��q����5e���c<3�����-ؠ1p��9��;�W^3�d�%B�y����O���|�s��'[L�������K�;���B._3t����W���L��m������I���@���z�v�6vL\pL���4�p'Jba�N�,�	\شN��Z&�~L>>�wB�������Q?1p���|�0=0������bA6�G�l���4���:_�G����5����50j��ї�n̂tCչ����:�9�i��ɽ�㢴���o���=��_f7��^<�� P����ݻ>C&���Ƌ�'3��v�@F�Fl��#�1�w�ܰ�ԑ�ª$yHS5�ٔ1����]��\cr,�T�b�:���B�Sa#���q��9�>�~�jf	GR�%�z�d捝�X`1Z�]g�	��Xl��/r���5T�>M'���J��#Ꙋ�6z�o<~N���ÉAu��TЄէ����F��2�N�VTTϘ�Os�`�A|�(���������h��r����b��dOfDx���_���ߍ	���C�f�@UT��sz��4�@��:u~��ٍVP������*;G�� �6��\���W4�ɦ�.ŷE%��������z]Ogޅ��#)������uKN$bY��ـ
/�f4�}/��|�Y���l4���˟TL��uV�6?$:d�#m�� �9v�-�6=�q�+�wZ�C%S%�.c�ϊ�I�բ7n�!�J�=���� �٦c��M��o6I'V-��'�t=6��e�{hPI���#4N�|1O7�߶E��l�m��nWΡ���{İm��Ѱ��q��ӝ����[��s��U��B$c��Tk�"F���s�`�'�!2�4�@��m{S�B[�1�%�Ń�p�U�d�bL!��@�e
,�Z��4R���u3Ζ�:�l�x+1 �5�wN߾�k��?����޽g�����րl?�n m�~j]�n,7�:.�������m��KTMظW����|�2:���.�fM7��@6�Y�i�%0m;��ZW3x�~x��1G�̽�e-&%K:w0�*�Nԍ����j	����k��k��V_�ț	(���W���Ze&}d��'Ϊ����au0�g6jQ�I�:R�#����	�6������A�C�5Ƞ&I���|���;�o�D1&�@�@�����1�T`p'Ǥs�m�����y���|�,-�i��]W�Vك.�1Uc���;P۪��+|P+�/�n4?�1Y5�jC˪��]�3|���(�CP�i޸��g�m*:V���M1.{U}�_>aA#�<��6�s�+J��!�x�{�܈�BI?n�O���R�M��� ���7�fe�����n�c�G���͘ODU��;�c��Y�:���� *<:�SK�(e�@���YE^�w&�.U�C�~��Ƣ�T��=����|��x�&L��< ��L��>ĝO
�rord$2#���r��4).�y�c	"�lSz�"��9�Eڿ��a�f}K2�����|]�9x��yc�����P��!*�,�4�l� 
��kils����}�&���H�g�m�	�i��:����щ�'�jPəa�p�N���?�K~�KM��FQh�t �i(�*<���u]����}/Pɣ���"w���"|��'�N1�����v�~�4�����75�NA�0���xSM���4�?�t���T�\F� ����A�"3C䓜�O3�`*U"���� ���+��K�D�D�	�*��/��P��%W|�%��C��+
Gi����Bb�8o�L~M�+y
i�(X�CZ@�.$�V����[jO�.�x��JT���f��u��z����U�a^$�tw��7k�&�,�[|qdl�[��b�������z7��ֽ�s{�X�6�It��E���~k��i}�����)Ds3ټy~?��(���du6�A$iڸJQgI�ɬ@.λG�Wï��S��د��O�$��r��
Ԁ:E�i ҡ�^.�b�u]�`/6v�<�a�7���T�z|�M�e������M~��E��;~�(��)��&��_[F`�6䔭`����X^Up@��	
-ɎQ��T�w�c�����b����;�:��n���mR�Hl�nE����L�AϳWN�����ŻP8Q2@Ǧ�ߨ���}����w�v=?k� ����\�ԶK����R�[��kFD�[ʯ��L)�[�J���+&�����E��Ch-_I�򰛒,P�pU-��i�I�$�%Q�(����:TV��`�Q.R����4��j���X"~����E2�rs��Ž7?���Xk�O�>P�ք+/���A����+������9�"��"+�r�1�(Uw����[5T�����&]�Ĳ���y�xXܴ^Z�ؐ�H�%g�>������x����-�	�2@���D7�Z�\�YЗ,Gk.� +�^I�\MDܿX�M���]�?G����qbW����sn�����f����t8���+�!��nV�Ҁ	i5�|����J�M�C�;➹j��j�!*��'-�z��9G�����������b�[ϸ$8�v��[Ԍ��cud'K������ap���Omޢ�.[ގ�~��o��&"��� φ�sȞyIHRy��V��@;��Gʭ��Ћs+��������{�����u8�"�A��j*m���Y�����ܐ|-��(>S�t&��U;�	j��f�@f���j�>�6MP��/���9��&���k]��<ؓz2���Rs���p5�dQ
K���Y�w�ѿ��0��AM��؄��V��ng �{�䘹θ�1��D^�iwg���ִŃ�K�\1�P �Go�F_��r(]	\��W6��y'��1�3�+Ms�Z�Oa3��z�_£��fl�-��1����%Z^�h�˘��C$������ڳ�p�	\}��Lpa1��T�ZM���*j��������8]R�{��)�b� ��oq��'����hjipx��C��I[�ؕ07�����֊S�A���_X���2#���'x��%'7��3��v$�A���َ3�p<3�s���{�;%����,���J�i�7����2�K������=8}r��0l������Q��6|#��Û��p9�>Po}�Q��.�5A
����
>�N2T<���w�4�V�ڠ>Ow]f��o�Gbh�4e6��uڈ(�� ��t�a��[�6/*:��m�e��F
��2��
`Q�y��R�Lq�5W$���h̓�º���Pe����o���rf���E`q��zx(=L"�1���8������d�
S��N��+�\�1�)B�/a����A=gq�%�6�����ӽ��{��{ף��9@ٳx�Wh  q������#j>����-�*v����m�^m��P�A�.'�<��,��^o����ݣn}i�ث�A{��k�?{q&Gi��A�_���|���T��n��h�!���F�\��Ȕ��*NR�v���𕊒����F#�+=A�In��Q�i�yCx%�J7�N���v���cL�)���F��(hx�z!��R�O��8���UFD5-u����ćK�����?&�)o�?���XV�L�&W��Q��]\yV���A�ϥSj�Z���]�A-����}^�!K��Q�V����G�drRe�����T	����2�3�h2��mM�"�F E �W/B���~��1*�N������\�S�9��Hu=<*J���ߕ+?E���Ť�d_zj,����\ў�X��kav�� �!QZ��t$%
���$��<?����%�ן���M̾k9B�	d���便��<3��i܁�����ok�uٻ(�o-��O��k裚G����w����5�~F����V�\�a�Qp��l̎w�t�R��9���D����5�:EN��P=-�Ld����.�AjC6TB����^�}*-iM=���$p������ֿ"

�g�E�:��/`�vR���&��(f���-�[Q��,g���3������[¬6���tb3���:�1�ַ��Ls��㾝����(bd�q�!�W��'�	��uYk��u�G�ꣁ0��)��M�RP� U��������1�X�������X+y'�g��2�� H.��V�QF�قZ%�k>�*
��j���?F�<�m���{� �sSB�K�����!R�.d�!�pz�L�˘���۝�X��@$Q���n�9������
�����2�o"ݽ������'�l�^�5�\�[�+��<���O�i��M���ͦ�I�(�g-��q@/4�}��x���ʾ�`�d�V3��{<���!�'�����1��v^�і��\E0��J��nUz�'Zsy��?��nLfz���"3�8��2&z�߲���}"��q
��>�;���m�iKꩱ�]�	�>�Dy�������G��a��1]�yX6�����!�ŀ.�6��g^*_�i�X�EV-�a}�V�`[��m���8��D|�/��p�}�"4�i~ݵ#<v#C�(�e���3���p�5͡<�I)���ޏ�nK�S��\x�PU,ex�R�~���鷚H89;ڬ�`�R�<����qC�/Pl��$�gi�h}�m�r���l�S�t�&\v�O�c0�爿�@v��f}#�ӕ�8_�=4������?�~�9���(�f2[��.KHK� �^�v��з�A8����P�n,�0��;�J�F�E��.}��,4�z�f�`
�n��Y��C�m�5�猎dA�y�>Ό@K��>Kn�|���}(\}�&@����*��i�>��֠�1��d3Ij$�;�Vċ����:�(�uao�SN�^3�k�	y}ژ~C� ۞�}�^����!i�诇��� m 3�j>�����4#gEY�đ�Q{c=`&�F�����EUb�t_�R*���{�.rnx������R����xv<G��^1�`Z*�������wnƼt��#��Y0|f�]�uU;:���eȸ�!b[� ek�#��6$	�
���1B�9�"����Ex���E7��Y4�b�����H�X�F�8�?��*R��/�g8���)N����<�z�����A�0��ϫho�Da��Ͻ�aI&-��.�/���E��ŢxHq���W^�іa@��m�F��6�)���S�G�:pD�O�o2M5}3c��p	A��$e��J=���崯-h��v����ӑqEl	�%�'^�φ��Bx��կ��&֡�)����Y�ɏiw�tW��0��.Ur�K�c���9�qYٟ��c�=MZ�迌/�?֣>���Z]C��8>�z�P�c�ӗA����&`kyĦ�k��A���ʮ梈�m�{8Jld��<Oo������pV=G��s�y4	W�"��Y}�q3����ypWϽ���n�+�^�g����qh��T���$���$�PK��g���kN�P��_3����� �lRBY���$ګ)��Q�ʸP�Z5��QOuf��
_U��>Ʒ���s�5�AyM+{*2��|��'�I��ʿ�5�����>��Z Z�@��p��%�z9<Vl ����.�ol��abb���㻧���gjԝ0B��^@,���.X��Z��Oh
��n��X�uzS]G^S�	]:�ͅ+���e@����H�e�|f}&6�I�l�
�?�<"��:�ѩ�Z���Է�m`�e���C$d�,fr/�2;���U.4��VKU'�{к��
)���/V�N�4~�<*�!	]J���-������YnS�0����ٮ5��[�A��?� ��ׇ1�~ai�1�63V���#��G`����h�Qs3E�JN㌉�{,NߨKR�F���n�A܅�{ᳪ�Y��}w���Hbv����#�ԎtQ6^
�/h�
�2���LY�'JM�T�M��_,t�\�gSvc�z!��Z*�с�s��텱�W���_��?R@��2����_8X_6\����7�)�C�qs��Р�֍.�HC�h���(}���Q�"2$<��v���PD���9��X�=���=0\V�jdE���������'@m������H�-ڐ�7	��,58��ڗ �:#]�<�n����r�	}�T�� �� �Ũ��+��6�#\��f��2�����d��zCjo��b�^e�i��Tw����W�+|c�{�{��{�h���b{�\���A��動�㋣�-T�w> Zє�ӀY��(�Or5�
4�$d���xى���h��Z��{~
ç��v/D�$ ���ʩ�%E��a��MB�B�����]k��3^��T�󠱽���1��n���ZS�ɶ�����M̰Drj����$�g�0����Z�L�,%���~�ev�r�O����H�eI॓e҇L0�Ļ��x�(���4�:�ܔ0\�������_|L-n� �^�T� 
y���N^+����Ć��*�\)���h�2�u⏡��|��M�'[��N^^�mJ�r�asR@O�lo#߳6���u���k��12�U�&���(�O�g,���Ɲ�T
�e*�n�yS����HL�j�,�,Ao�q����[{�+�<޵A�[j���W�F�|ѻ��`���'��]��'�I�f
Ѩ1����浚!�&�?.R�~7��6�������y<+nKhD��߲�T�_v�0����IY�D����_T&,�bE�)�#�$F��w߯
�^��͢��	�&��)T���{�����v�&_Ƽ�Bk�Un���y��2#C��9=F��k��0�E; (��_��!��x9����^9����c���"��i�{+��t(���S��@)����9f�꘭�,�/N�Ӆ�E	�'�K�%:>b��$�V���Vh�E�d�l0��c������/d�;��[�W�{4S�C�VTb/�9 ��S&��D��K�R�PU�����X_����������\�,����l����ҟ�	Ju���_G����<ȼ�����$$�3�y9$�������6�;�z	=�<�;�����ޅnV��M���^�vXR�Ul$�.,�hR�Ԫ��r�[�t1W��/�p�&^��U]U��:kUu����="tBt0p��uf4H�G��L3�&�y:j��x9����Yk���5�R2��u�1.$���C�G�����H�cR�E�1`K�P+�צ�����Q�U\U��^��g{�t	���2�.k�}p̱����@�w�Q
����'~Ӷ0..��B�Ⱥ�m�<eP�:�~=���R�T�3>#��˘���5�-�5G�q)ɓ�|&Y�:@��Tr�
cgn��$]8�����`jm9�듶�_����t������-��@n6Ƽ����ğ�44!�=�� ��!o]��4���Ѐ��m6�Nj)RUAT>��M~�N���	����R8p�N�WP��[�T���3.s�U�+٨���)�o	^�;�HF���(���oxyc��+}��U`K��:޴·�rqJ����-^Ns���7�K��l(��p���1�6<��w�HmHD�)R�d���8~�K]?�8�j�KL(��x2��?"���f��@�N=u�͡�m�A_��z �8�!��}>GA����+���m�|"ʼ�������`8Μ+}V�{�ve�w�J �/�u���7״��h�~~�NZ�W����	�����ǔ��t<�A�j�kEmq/�rg�櫇E�t�Ex��ga$��L'��ʀ�i��;q��t[iy�{��,<�MDJ�Ig}��]4T*��o�O�;_���6�����'@�B��[����0��Z�c+7X��g�"��r{0g�%��%Z���\-P��i[���f�z��k��['^�h����z�������ܑ����W8�$�v5��~L�&-CK�kh+Ȉ�i>B�3ŀ��v��+�5���H.O6Q� �
f5D|͓������B��P����ՠF���!7��Y�8ҽi��9��kGhE��;)�v��_ۚ�gl;�~�l K|@�kK�"���0�@(��?��->Qftx7}�Rc�F4�^s�L6��c�??��nn5nh�e�$Z��N�zp	�vz�fQ�)�f}i3��������
pr�]��k>D��[l�{	e7����dX�gY�
����4��6�V��&܍�p��4ԝ��̺�"��>��Q�+vZ����OlJR.��LnMj#9�US�W?��2��V&��*�Ow�f�:��)�!ǋ��$��u�}��+�zڤN6�l�9�
J��6و��Q�[�l��o'��K��4v�ȕ���=�ǒf�/�xJX���$����_A�▇y@��Gr�[16�3ɸIޖ����ƶ{����pT!'��@uFn+�ӋW�E�Z��~���M�{R6�ڟXI}Χ�NI�i$���]Md6ؓT��h��0b8�cQ	�&�����֙��
���!�	�m&�b��/Y*����92S\~�1�5$\��q�W���ݡ�y���n�O��&��P�9���q���GO�T�Wc��[�j��ܰW�I7;��(К�ɮQ�t�vh�N�	���z�*�>�^1Q�z(	}{h��.�:��gE��i�$*�1��L��Y]�h�J�aנ�Nw�M������ɪ0�ܚ����w�>�ZH��]A�ޱ�1�(��+~|���d�q9��*�^�>�Q�z�_1;�
�&���n��g��F�.q(3mj����Ð��Jx����Wi��D~�b��u�^O�8jU�N�U�%1�<�����~��駩p�@��V]�0�d7M
�z	��<��o�����~p��G$?������T��z���si�v�m8�~8_ŧ�Bg�������n8�]��k�'&~����V����o�*Vx��Ǚ�=b�J�$�'�2͘�� w�d�]Z��!��Q�u�Yi��;ǣ�4|��6=^yQkⷲl�c���ގ�K�>���O.�۽k>�xDO�,Ȫ�����vߛ'�%+2#�密��	}n��������L����$98�����$�̆��󳾔dF����9mS�M/����mbf`�b��C`�N��x����r<�D��kp>4�����
���}�΍q�����^�G����n�� 6��hz��y[�}��-��^_f�z: ҡ����M6�R80��8醜�V�*݃�Pgۈv����<'����1�[<� ;�9�1��˕c�&3$7j�Ϩ�|���s�`_�|x��DucX$����{��G�V�pG��*�¿[ս�[�}0��4ſd�X���94b��S�t�ץ�2 � ^J:�*t.z�+�%��
α~ɘ�ĵn�b�
s�.H�vt�XO�00Y�k���W�i�"`	�d)5�u�	4	�4졷� �!+��e=�L!��U��?8d��1Y.��e���;�M@t�5�(�õ���d��u���_P���"<�.�&���:X��=�2��e��f�>�n�����;z�
z�2�&�L
�7��e���jD�^�K#7����t@ �R����Bȿ�f<����Y�)�mŘq9(fG��fa���|<͐���;���(H��6�)�����fT9/���5�W�6�5{��]���PEe�p����9N��v�������C��)T0z���)�N��_�����j��a@[p��
�
%�0yOﾬ�k�w;*�^/�y.�i�L�Ro���hZ��:&b>����<d�<�%�	n�He->D�j� �\�Hgb��eEZ�Wl h���u�PAJ�}��H��]��?ϛnpW�]��ȡC��*D7�Z��'8��8�Մ�E�u��P�Ǻ<���li?�a��)ـ�%&�;�BG�)���:��,	���c��L:��2�T��E������1���Ef��02��3���G�)�g�c;�9�V�� ���ɿf�n�����'9x�^	>(ة�}�h�����yW���1$3z:��\�α;�Z.&44J�U�%�qb�u2l��;�1���󂞥g�J@.��ns!5�`3�ē�p�0����vl���<(�+�Yn-��6O}&�NJ����,��Go�e����D��N��߀x�Al`�W�Vq�����a����_�g���b)��F�T�t�⟌�Q��[��t��Y�D\�Yvy�.��|5������΄����+����.�c�e�8�jS�ZPM�fP^3�=vd͊j꘨������;:p,r�IL_k6����ơv��W*��EA�(Q+Dd�Ǽ5�Q��/�X�wc��ﭗ����8�D9I���	�-9o���v�%����P�"V�/�_�Y�[7[3)�J�@�a,t�}i:���2�5U6<@��Kn0�;��,▝:Žh�B�x�]��kꯗ����=[�ysaK��\�06cH�;ȇFJΩ����~E��o4=]��Ɩ��>��Va�h��ٰ3أ�],�Y���a���}�)5A�H��Pewѣ��lQ�d��=)�/�ny�
�(^G�D��N�:�6�uȎ���+�f��>�{���
���Q��}��X�_)^��_2(�~y�^�	����^�V���fG�R��}�]��ܪ|�����hW�Zr�S�_�M�j[?�E��٘[�OG�N�2��i�0 4.���}�����B�bO8z";x�&�R��ӯO�1��>=LVȀ>�PG��ㄌ�҆�� �VW [˧�_z�
�Kd�|����3�	��i�_Ι0<]�Kұ.r=؇}�K{"˸�
��Y�M�#"�|�����͒7��u[�;Z̑:�5Y:�>G��ѻ��w���I��<i���f��#�S���@��ȣ��HS��4�NBͿ���/�d'Äƽ�l%(��Y��Y��\�O�N�:^I��ɗ����
aWS�����Y����rw!�,\mJA%��1]�@9�ֽ\[��bĿ'Ld%��<׆��<#���!��V��d���-ɨӐ�f)��ҏ/(	t�K�A�?���vVr���f��_�+f�����$"�>sa���j��c.��yK_Lޠ�]Ek�c��mK(��C�}�$�c���ܮ�e�xj���������䤚:vA?�֮a��-2�ÝB��7��G�㟃Uz�>Ʒ�KLE���1O�����l~�LW�Ty�2���>�6OL��FU�2
�(����X�K��~�('���Xs-6�QFY�D��g�̘(#IA��Z�<����0�>!JɆj6�'�s*(W�"H�ƕi$��wB����B�-O�§��ĚLl/��.CC�~x�k^�ºI�ͧlR{��w�X��~���E�.e"[�yԉ�%(�F�~i|Q?���4m��0��x�΀M��ͳz��D�Iq�T4E��(����Q����[{p'n"�W��2�o�eEkv�0�.��0��_�н�%�4S��.򻆊T8*
�m�V�>1I���,�s� �pi�[���� �%�Ӷ����s���L3nW��LP���L*xh�AB��r���k�t,��oO{�?	ɯ�1qv#���6n�� F���b�+��N\����B�8)��0#�=�.70��6Q��{��#��d��+
��Cc�F������ص�������em):�)���5ځ�Iv(y���AWb��E|t�B��A	z��mp"��h�o	���SJ��A��
I~��L�+�
n,�u�㰠i'�	��Q(����|�%.*/��KՅ�^7d����E�9�^~FlA�o��k�!/)�	A'fe�·���+���y�7��Bp�h>�s9��m��U�1�[���Ce�[k�����l��1u�S+;�@CJ;�t0n�"�A5��%��>�D[X6VS�����	���PrlK@0^kJs�w[�i�MLD�<��gy�I�� ���?!���]�W̼�wg
�±/�J2�D&��*n��Ɏ;��bHb�А-8ݘ�+�ʦ�8���\>;��c��q�`��������&?r���Z��V�}C�e���_��_fl�:�Ё�\9�
��D�`}�ގhA��� FS�C��F��w(��xL���@��Ӟ�0�S ;\fQay�<�G.ދ�}�s֬������4�ָ�6^�go����<�C@���o{��`���%bH��{��.��ߦ�T8,�͖�Al��%�,�In@�Ө�*��BC�R�!�a�X�S��_5/��l��&\��J�/������Ǭ�N�~���յIy6��7��
�XEx�����`�$�M���?��йv��Kd�c�o�-U�\{� >��}����~ͣ&(C���YW"4�<�I��"�P�gã���j_a�"�/yQ&Iٳr���E��c�ԪId�̘Lᬔ?���g�H��kroNmI>z�'�q���:�a���nmH�����rl�(�3��!Ekp@��0�s�_�F^(P�?�(0>�i�i�
�	�5�W�ݮ�a���c�HduI�?��z�sXD�d�i�ș`��7�����\tU]�(|����1�v�λ���#z��i����2u��(j��]����#O��ˢ9�fǧKy� 8l�M��"A�[p0��Z��R��P�Q�i�9�%d��D�KYy%E����|lE`F�H֗p�z%��� ���O/$*���\��<p�Y�Z��NÚW�G��'�"���[��I�UTt�a0���rx��M��
G>�㨫����VP���d'�0�e'�G�H�z�oxA�QL�G�Jn����Ɓ�|W���E�۪� ���3
X�Ƿ�����4~�&p������ࢽ��Tn�mD��.:y�o���7ӏ� ӭ S��}�3�i���i�Y1s;��3�V�8b�`�s���!��Q?�nK"v��o��9�<�Ki�9�#{��ҤD�L��w���1:2BJ�I:��� ���~'��B�	-�L(��nrX�%�^����BTas���e]Ay�9�����%ē�E.v��Y���"ȉ�;o�#`�
U���%g���
=5cT�������?w����4���dM������9�y8���V/�u��焅O���2aw� ���H;��5I��4�ק�O�])P�@��(� ��>�&��db�M:R�yg/n�:o�`'c����Յ��m�u��������33�b�Z��n������Á=`[�8���6�F���~�Hk�_1�2��r���Ⴠ�nq=��^z/+�ĥ �Y|��T�o������B�{.*58��|Yt-�@b���A!�n��M�J��q�rk��,������0�#��T��R>e�V�I٥�=����f'	`�>۬��Q�^>Jf(8S��+*7��E+h�X���ՅY:o#~�$ٿ���
s<o�����@�5�xm{�t&����ףv��C�J�~���� ���6�L;�� �O�q�H�Pɕܖ���<(�!ޡ��j�h����<k��`!
�44�4MK`/O���X'�ch�[h�N��f=gV"��_���8�=�n��1x�k����=�S`_+�\x
+ Iҧz�t��$y�&9���6i�#�gF>�5p��{ƈ� 
I{9{�w&�|���X�̊����i�V���:~��H�YO�&t�����9#-����co�\yYs��䣉�J������v�
��Z`�H��>���8l�+(�m��/�#�?���鶷,S�%��p��,�v ��y/[�QI�n0�P=��he�P�jY�z�<��M��|��lnP>�0v�W�tENR�6hR�<^���4<�d�r�k�d쇦LhEtF�Ӓ�Ј~���U����f�jN4~j�g`�:%�ㆁbV��sb�L�
'{��6Tg��j8��u�_�3��[�炆�X��훚�.j�Z�a3��,�>��wN�,�/3���ݷ����i�YZ�`Ƃ^��4e�?*��)�K�3�bI!
�x6�2(цQ���z~����(?sf�ڢ�����z��c�����I�`���aQ�)ehǲ�F.W.>�6��)np��Y�yP]m/F� 	��bTaF|:|�1.A����H�le>�+�I���)�pp�'l�׮ڐ���z1���u�/����wek3��e4�ʜ�Q�H":3oo�ְqU5�vUs*��]a}�Q��q�f+�Ma�}ۆnuW�ǅS�o�p(�<E[;�:B@�C�/�fq��'-�g���,���a+��)*�6�P����}RύRT�����REҨX��}2������e+c�O!�4���k�{�Q�E �[�u���t�c+�����闙�h��{4��Wy%:2(IE�7�Ѯ�ў�{�iu�Zz�m�$|"}�H�?����Ԝ�������t'���%w^��b �N������ko�ZX��GQz�R��Y��z����sA>��J:�ŷ(�^��DG�A��I��S@ȶ��,1P�)�UX�O��}s�ƿ�#\Y[�1]:<��������@��  xks�L�4	��-�ނ�y��&?��+���ML`"Yޛ%�l��j���Kyٝ�W�9v�s�&H.z�k3����G���҇�:�Uel�^n��W�"���>בY�acuC~8�2@�e{���0<W�X��*	����;��C��*������pQf�?�1"���r�uŚS!I���މ~���DT�b�2��U��_ITE��<�hr^`�0.��2��r:'ժJ��v��c�h����:�������}e^%�]��7B�^�+�v���10��|D�Ga$Vr�O>�<>���D*>��I��5�
�;@DL�L���i@�r�=��Y	0��Q�g�Y��<"���ꟂW5Dt;UaG�њ�Ea2F~*#?�t�K��(5��yL�W*h�_�)8��.��h_2��'�v�T�����n��+t��AQ�VX��[׽�6w���Y�j�(���+3��37�M\�m�I�7����`|���������ȼI������5�gE�sjG���t+Ȉ���(���*���^���������[��3��R��M�E���r/���ᫎǽ����^��܈��-ſ�X�&�d������`�:´�XD�7��E�� R�P2_A�L�0��P�3�F>�T �I$b���q|�t����~�f���:�����BRm��)�6v�����ݚ53��MJ�	鷜l��?�@L�gn�K��k��v�h�]��q3ʺf�t�C&7:|�Վ�6���7�6�o�B�8��7c�P����%�?3O&x~�;M��.8Zz%A2�ˁ��M��&L��z�"]X�<�
�o�P�Ai{�w	����+eޠʽ���2_慀}�GL�u�v�y�	���a� �9�E�|����g�f;���P�h��<�JR��m*/P)2�۠��m�\p��if�󫃸tf�	��������B��^"99��2��s;o���(�?3qP��NѬ�oџ���]����*A�=I�(N�����rc>��Q �+$	e�}�*����]�u:ީ.�����Rtɔ�:c��������*v����N�F=� R��;�Y�mz ��. '[35f᬴�N��޸܇���?�t� �bC:�?i��l8��,r��S�tHG؁-50l����*R�m�z�^HU�_������ 4xfrd>��/Z(���by�C6�4�|J��Ԇ �U��D�i�]b'C�vd��kY��XO� ��\.����iӝX�2���.v���<E�6}
��zp"J�1�{7,ޘ|݃���6w�G��Ç���N��]d�V�((�R��l��v�Xig��ڪ�vQ�m�b�=
�p1/Q+)h�ڂ�?$v��&�Q��\�X��y.{M�:���Wz[Op4/>��난R+p�Z�M��p(�/�o�e��6����2d��;����.E�.ћֳ��1_��dp}���L��v	U�6�1�7d����9��\�Mo���K�D�2���b�yS}|�A�OJ��s����F�A���x�*D��	Ď]>+�ʚbX|� ��vH �X:�:�qe}ʂ��sK�psRoΊZD�ކ�b�����v��X��p̌ٗ�H�Y���R6��j_dh3�
W[�gW�J�#����\?@��t��[ JZ?&ɵ1���B���������5�&m6���1�!�S�s36K��*�����73�pqUQ.�ZjR7����sq;�3,ϐ�?����2�� ��~@x w��C�J>����O�]���-��5���qC?값��}��֓��|�ŋ�1��d}NO<a��\�Z�i���R4�&6T`5ض��wNN�E�]�����[�w{G��^����Dѽ|��\�Gfܾʲ�U��yĄ�2��hzL�R��9I�i������+����dl�L���.O��Bշ+�	������=�22=G$�(�~�p34f5���<ӛ,O���hv��6`6��S_��%��S��D�a��*��z��/�J��ۅ���3;\5��'�����tJGa&E������G~�S~C�1̑)��MPUO��*�����	P ~�U<��0�A�!	�Q�T�Wn�"R̕,h� ���l�BK
�_3H��+L����X�N��AN�~7ݗ��  ,�����I6c��K����MAi��$����M�!�ҋ��0/CU�[�>4�ό�=�VO3��<��7X�G��1�#Lר�NXF{�1���{�� c�^�4�-���U�L���(`i5�۫���NR�eQƁِ��yP�-ء�_+ڲ�E<E@3���V�퉶:�J̺��z�/bz쩶���?��Χx
|�v��@�>f�ݗ	H+ZJ75^���<�/nӰ%�WdK���|�����U�q¦�� ���S����__��γ�K���+Z��`�F��K@a�)/���e�cX��@<�+OH	�����}�P���+a��+��a�dcj�m7Cx�㱳t0oEm����:#�����/Z����d�@5����P#rJ�px��|ӆ�1����l�m��9�O�r�1�x�m�7�(�%�K\#z;�+>�����ȅ����kXCdU��J�ms�x̑Qݭ�t��>`H�5�T���j ��ļ�Tod�}�˚l���.����_&��N�q�l�������P�P%�]�;��Vu�S�c6���B�'�)t�7�:
ǲ�6t`��%��I1y�-B��.c��F��2Z�M0��(<)e��'��xgW���\њm�.ě7z�vܭ|C�q��Es	�i��ؒ��{G=��<� � D?lB~��+s��V�Cy܏G�~�/|���pl^O{\���i��Ϥkx2OB�K@5cyx�2�p�=�Z̑j�4}t���H�?:�ko�
�r�����S��~���<zJ�Mhy6:cfu�%�]��hۊ1=|02Qg~���6__�\{u�P4���x�}��S�R��^ws2I�QZ���/���y�=#���
������k�c��,\@���L�ñ�h�@�U��ޠa�ƅ0�I��O�c��a����,R��I��o�Xw���# cD��Dؽ����g��ޝ��E�<��t٢�����_�LLQq/����!C�͖c�iA8ߠְ�jZ�U>o�A��*ǠP[�W'�W����&eB�fp�!Y�|�U���.cHq��K�
XP}��Ӥ�IgSD��
�?��r�K����)�w��)O:r{"���7��C9|-4���Z�������՘�w��[ ��ڮԓ9�Ɣ=��	E���8�]M�iv�����|&|T:�:Z�$ �T:aI�%� <�uv����L3u)6�g��	���@DQ��5���R�t�x�����"��n8�T`�9NB�%��u�� s�-s����*:Ê��M�8�F؀&#�&�"&��5É�K��oMd�҃u�řU)5K�s������Z{�(&9�3�{�b���a�[�8�)������y/6�тkg-�#����l@ȷ+�����x/�LNY��x*NZb_�ƀ-�^B/ӧ�>q��(h�x���d"d�1ǭ��з.�5'v$MJd���Ac���� V������||	�>V'��^Ϳ6�hz2�3��@
�:R��pA
vOt��A5�7M!z-�X!���KW�����80ب�;-�Q
��4~I.��i)�@+�N���������T<���?�#���d��6��bi_t���)	�ΐ�%��L��	Y��:�@�o�3�HZU�<B����e,1\��7o�N�3?t�������3.J!P+����Շ�%��x�j����X5�!�}#�h�8{�G��DJ�v�{c�0���:Z�J ����|�.�D�'w:¤��B
�K�V��ָ�j��z7p�r���_���
��")��>.����jg�9%��
&�bȅ�Lr��m���9΍�S�A��PE8R:K��ض<�gH�H�f�~=J�-�Nѭ[����|հ��MlG�l�ƚ�xJ�u���i���
���~�i�t�s��� ��PH3�Q,sL.��S��˂b%�� 5Gɿd�1d�X&'7o�>:\�X+�!�蕦����ƪo	6Jm]�?q�G�3�f�w�n�N���%�15��*=�ܤ�b�p���ɉ�Ɂ�p'e9�g=�?�f/�E���~��u�w�ȓ��qI*�|��Z|�`������/x�2>�C��\^v۔�~�.��Q��x�l�#22X;2/
���x��I�M��S�̻ۦ���î}׍�/�[+O.-�3�g�1���DJA\���P[���m��9N}����G�Ao�0e߷��C���	�El�6,KO<VYm���0���̳�y����)ݡT�u���+�Ƭbc��/A>�v���߄�܏ ���X�f��7̕|Nb|��e�"P\�A%g�дn��P��L��)�x�U�����?O�2`V���̔�֞��d1`h��� H�Ї~Ty?X��3<��)T؜��Ěî�7�OF�q�tn�$ᇟĶg_���|���`?qs�ǭ+�H�6��d�Ϭ����9��(�H�1"�70i��$k���֟l� ��u�+�����k���X��6����%w�#�8GvE���9� ��d�b=���q�א�oH4�R�@�{l���'�Òk�� ݗ�������z�sth
o��t0+U��+��Sq03��Nb���?)��Os�W�4s =��pX�cNA��.�!�HRC�T��uT�#OP����+*�5�.B�xdS�Neg���f
�ؘkO��a��� ɳ���V�F
B�l.����o�dȼ	�m=v�%�M*b >O�EɹƦ�Ta�B
M)�`��iMV�>�y�Bo�@�yF�9?)aB������o� ᫯�8Qb�>b��p��{�f��5��z�SS�bJ��J�%c��ѵ�pqL9��iP�EA�wA�[�U���q�<Q<J՚�F��(�V( RR���!��m➚�2�ճ�vCf��(-K�.�	�K� ]T�X���;�k'��0�ݵ�e��R���<�(��t�"�}��ț_B7c5q�Y��p1x�'8�b�J��l�8��3b����  y`����D��>����/�^~�rv�sy�
�9���BA��0U��%oY��xWB_�FXMa���5��B�%�Y��G�z�=�<A��/@�e��/�v���30�ҖN}�n����/@g���#�/����e<,j�:�1���hhux/�X�h�f��{ŜG����QB���g���e�I6���]�0m[9���@Ҳ�uo�s�O�������;���
����u�Ӗ�A� ��U|��������Ϸ�}_�����nZ\��;��?�ܘoV�8���l
�du�`��S!����b&P��r�8I�f�7M��E����v����y�@�UeA��:?.Y�����FB�UK_�"^�k�d3Q�8���}�6(x۠9L1:Qf��0����ܭ+��W
�7��R_�}�"��2�\Q	4#1e�<[z��XZ&o&�b����71�mLt�<�����妕�r������>��iL��@�a���I:n�Q���Jlr9|� I2�"��,mL��ψ�ٮs2lْ� Rݒ $�8黪گSK�Rl|s�Ks*ԇ�4��xP�PN^U�D�,}n��VMssZ��;9K�wZXv&~4���vv�lϧA��y?����{�y�I��p���{IW�G��J��N���+������?��0�՘�,s�]����'�YH���Nһu�ܞ�a]��ze���B7x�ŷ�ӏ����aV$�������|��m���o�d�̕�����ٗ$^(f� ���21���l�N���l4��s�M�F�& !�IH(��yn{�?q�ݜ{mQ�`�j;�T=g0�Ћ[�y�B���� 9{`��6q�meh�#�����Չa�2� ?۫9���)%��n\���%�v+���ϙ�n�ɢ��6`-�׀��}��v���D_�^��9�7P�5�E+p
��LWO�]2%&DԵ�ݳI;$ٕ�Nj��� ����$ϖW�9a=�����a��o�o��7�f�#�쥦�!�?b>xz#5;�+��f��ۓ 	��A�.'�왬w�=���v�>��^@�H+a���y�5��䳻Kf�"��v+����W�e��'�$�2�(R�]�Y6��iktm���M�,E���A�6.���IϊH�7����y�L1��S"�R�>T��a��#$��h#zg&B{����:�H\���؝��W ꓦo�#9�TX���n(��s�M��6�s���Z�3R��.z$H�i$�qW��d$Zs�����3œ�ЌZ�j�hڷ����b���}�CH��+W��Qey�Be��3�����S%��Jk�}����$(�|�į��rpٴh�u1i\k}���ӄ�L_�;��fL'B�Z�$��Dc�\�n��O��aX�pp����U�;:����&������w����k*"��U� $�4�"���n�X�@[�=�Y�PV���Pl��	�T2+��C�"]�f)����g�5�zhJ���w1�20PS���-}0���v�.2V�U���ZK�5�z�j�Zl#4��$��2�Mj��,�"��"� ,�������J�zF'��wKV{W���*p�ڱ�1]~����U��*8,wJLB��C��<���V��׍o�t�yϬ��`간��`�
�c��_���(�o*�g:��F��h���֎}��M&�����^�i�����M�!Y��Z��Q2qN��^$�Հ��,]}�"!��i|mI����jp��Z�8��L�t�[�6j�q�#o��w�_2ne[8���Q5�F]��.�'�L6�o�ҧ�l�KKܛ��a �h�ё��xA��6Ḑ|�|wpᴚ��8�-��`�N�x���2`2��I�/�j��V���Q����s����g�xj� v����--�a�p���o�E������O{2�;�~'�籰ܻ����G��1������fI�Mb�Z�r�Lc͎�}����Fr��f#䖭~%�jh�/���C+�%�X�Y��c-��!�X^O�?2�����*d���U��ŒUM�1�6c��	����͑�b��K�,�//�!��ԙ��Zr1y���b��iΪ�1�K����;�(BZ�}�~9�"��W+�4���c�ܑ*��냍�m��Af����Gq�+I��*v�U �9�@����H}�K���^;�"+}ƨ��t�g������R��r7@�&������'��)�G@j�r�B.�v�]�Z7Bs�Z�O�4m�v�s����M�]�t+	_�O�����O��"u��}����/û)���p�m�K��q5��Fe�瀺|z�V��~�3�����4�9܆������r��h�\�|�#�qc��ij�:��F}��#���1�.*���K5��VvG����9��Бi��@;;_�
1���F��Y�;ť'�`���V۬�����i�q$�׻�n�_��/g#�D�%�������M�/�V�T��'��_T_[������?�� * ���R�x*P��ߴ^�0`��{E��G�ѿ�V�wLM<���x�v9��Viz�he6��+�b����(���y�F�����:;�L=��l��{޽��h_��Xo]�e׏di��.V8�b����Zb�\�{�8�&"���Nw�1O�N����C	�D�M\fG��0.��y��"$_�[�J�gp�qp<���<�}D���;�a2�hmo�?�o�Թb���N�EK�ҋ7��Y�k�Ǟͽ�(;.��A���T���E�lb;
7]�\��3m�1S@"��o����}(7�P��L�D����+]�M��S����n8�n� �G`���׳0v�e��	���+B���{�|�E*�X�u4H�x<�˪Bx�R�{�H����+�i$F��09+~=��W<���E�Z�)8�1Ya����ΠV�H��t���}����C�'�sT+�M�ֈ��D��B��u��ج#��[^��ۋ�B�?}6@�%oB���Rܣ���f�H)|��"����qn�j�ȡ(����L\��S�ퟒ畒F
R/[ltz^�� g>��sk��8E�9�1r.�~���%n��'0����9#=g�]XSo����nJ�;C-i:q�� ]`�[Z�ٛ�
����G����F8f��>V���V@;�� FPȽ3�N�� ���?<u�r�':[`��2Z�b�P�S��=ױ��n0FzB��L��k{6�,b֪!�-i��n�4�ɣl�;�,�1���m2h���P�"="�����w�f�Qp�2{ŷ��gj:5�C�E �ƘX�����|���qB䇫�DX�LU�b���C��+�T�,���<�D��D�����-��X_I��|�P���>��Yߛ^��-T?��_�@�k��E㛿�4���M���D���x1�ݳ�i���N�3l|Z�1y���5[,zD����1��MPF��W�N��IsK�}z;c|�-�6Z�x]�\�0B.��h��.���k�U[7P�[!�{AG|��0�U��S�;0v��c� ��Ģ����a�[8Ъ��t�Ga�%�Y�w�9��]ƶz��W�zmR����輮�[17���E�
 [C��mi=�:�'�X{x/�q(��^����s0�� �]����^fb�U0#� >R�XK�� ��z�q�-m�8��O���3�e;��)<�ˊ�Ed�$�U�@��DW-f�\�+Z����;K�� /�.z����A�i;�+�{{ކ�-�8b�LS�0�s�O�qP�2w�
k,�*���g#�7���Dg�[M|�qzF1ʛ���f"�Z���Y�Rp<�a,v��*O�q����B ��Y]R`�Gd������{2;��"�չ{��P�$TwE~У-�����82���������� ��%&�\��O;� �~���j�DY�j�W!��qٔ��z\%?�2�&N�.�xڏ±^rRQ�ߨ%#~�?-!m��q�)b���	�f�9샬�8��������e���Z�}��Oȏ2�zr����l=K�巁����@d�K�4i�m_[=����t��5`�O�*u�@��ĝ��zؿ����
�u�Sg��߱�>q3�h��%fd�:��pJ����%ی�L,ڌi�*C�'!6)��"'R� ]���Nb�}?eS�# ��g(����xZ�*N�z��g�I���L_I�5���#9�;�
4�,,�	�#������H����(�%��jG�ml�DBʈ�8����ʣ�k���t����A���o��؂t��_� 
��l�iX.Ϡ�ڎ���}����^����,�ul\�[�P�P�nI���M�r�f[m1�.����6%W}ډ�]����\�����'��x{�S%��F��Q8��_��\U��xi|�F��y[
���h�9���46k<����zU�9�_
�~^���m�K�j��b��wv�0^����׍�1���0ڽ۔� �Z%��Ii�[`�CpF!��W��[D[f���׀�n��g|B.r�J�r���:
�����_-u _��g�0�� �8��Q�G��6����?3A����Tꫂl�����棛��VJ������+*��r����A%`�P�!-a}{�>zD��7�"]���z����I�~����&�7��Ҹh�O���L�AQD�W)�AN�Jz��!�"�ḷ�Ř�`9]��w^��͊)����}��qM�w���H��uܪ���i�i`\�j�lO����5��/�)��6���0��u2��y^���{�{���k�C�p�2��A���
����\�@�5�j����<���cX�>T]�j~�V\@1�N[ �/��W3J��s�_���_-_�DRT���R�$HD9�l�8PY�c�lE��������W]`��C�{#W���Gd�����T�����?��T�Ӹ��z�;��p`��{t�� �-&��S��(K-���vS�Ӡ���d�4����?eLc_�ZYReb6��ku\t�Zh���F����ӑ�<�n�3?�$fo&���n�չ���S�xHu�<� �5졊L�'<�c05�j��3�D��	���BnꝀɢ`,��O��oR+�/A��C�?���,J��]�V ���JAݑ@��N���/����u�{d�s-ī�D��a	i0s����it�͒�o���(Y�RZ'�<&���T�
F�W�Hhl��r.[��+/@�K{	�ؖcr�`���1 8N�J��Xq�b���.�q�[����_{3E�����\(� 	��kU��"�2�"�L�pO��T11'޾QƑ;~�JO�I��/�M��ѬD�oW�
]W�jk�5��3�I"�k�-Y�oc���.,fJL�@!�A͑�ѤL�������!����F���f���7�>���H�2�Z���B��>�@'����l(H<�U~]�}�,UcY�R �Ǵ3be�3-����M�����0��O���u/�fh.ZF���>q�b�T�*I��8T'|c�N'�\{�|Q������i�%^��[�ά@F��RCR��#��uVL�ñp]]��ُ]9�c,�
�r�c���������>�w�Y�𵿞����#&:ʑ6��8���Zr���_��M]|�H�V�S��qѴS�0��%[!:?�����M���Ҳ~��cZJ"����.ƈ�}h<b��Y��1�����k��J+n���KlK[��\b�c�P�����.6\�*+�d�ߏ���(��l��F_�"~�Gp�'b�7����d�������w��HD��8�LX�y,\�鏶�U��e�����l� �l����������4��6����K߯5��Y>�.�|��L�K����Oi�?i�H���m�%u�����r@g�+�Ʈ������0nd�{D|@J�4y���\ ���w�����[��ۇ�m��d�Dx�o�|�������$Y��`��
{���9vD��m(�=j�QY���> ��2S6�nr������a���u��+�A����V:�he��ҝ���)s�(N������p�����Bېg6�8Vf��aDC�lb3~zx����C�d�EXz��eU����RRЖ�1p�4�����TѤVq��^/܎n�h��4]<QcX5��Qx�0�5��_
�-3��Aﲲ�}agp/�Z��d���k�c�� @.a%�`Xj�Y'�vA� �])L��;xJ=�b,
�ƉN
��r$�#��g.�"ϮZ��h��Q+�:�-C�C�]2�*�i�T^O�2�J���d��;+Z"��3��f���9��n@V/Yϒy��U�ZD���}���/lű��&�3���Pkҿ?�v�>]py����9�fr)�9�V�,�O���u7_������7�/ ���������u�� zj�m�}+�Z#��Q< F�U�$�M-D��>૸1���JPN`*�!T&�v�y��}�#�tWf5�3�8�����1����D͟�#<K������`u{^-�dռ��oE=j��b��� �_��edL�����US.��RՑX�͎4Y�.���?����Q,�{[ҹ�k�3s�̨[��(�*߱B"��pĪQ�C��p�|�
?vP�d������n*�b�qJ��IL���h�M:��QF׍���D��<5�JTӫ%��h{�9�����s���������VU W(C	CTϙ0w�?�KQ�6a��cl�����dY�rw�+�E8%��O�'��p%�,����uV&�9�E��i�����t���=�ʙf3���Kf;�z�M�'@nʵ�I��ﶪ� ���P��uS�*��̡��k^>����������U�sf�\�|�����՗[��&�)�}Q�-+�x�������~Z�5Ĕ�(#�&�?�9`E^;��ym-��u&7��,��-9�t!�O'����������?ݳ[�El�H6"^��O�뎆l���f/R��� ����n]������К��ْ�����K�;�<Љ�<�����S�o�	���P%���?�\�}e��F��x9�aљ�c�D�~�H�	
�����49f��xk�]̰Դ,��HCa��Q#U	#4��?�mt�.+۝OF�jD-l�C.�J��:��x{�*��$�gv��ɢ/�Ѽ@�S�VٺqG��*���X8�O;�;G�h��e��e��UL\�'�>#*G���	�NKG!���ö[j��C�m�/��i$w�[�	X��i��^�Z��l ���R_g
���R�a��T_��Ee���=�+��&V���mdP����FƄ+	�}�s�����t���G����b��I�Cg�x�`��Ԥ2�����4���%CS{���/V,� �$\yt������}p�۾ߧC����Zj^�����e�6�xh�V����gu#��$�g�(@�����T<�\�Ֆ�z pT�>�$�K�C4@8�7]=����~#�Ӿ���^B��O�;뺼�x�W�k�J�q�9�1#v�R#��G9b`���k|[�|��)������a��a�)��.�񯇡��uՋ���V�'��yS�X
�B��{�6�H�_v��q
o��7܆j.]������.|G��l�p���3=�b����^�!>�B���@P@�)f���_
8���~dh*O�_�Ҧ���x������?��KF��M�i}���o��*���*�DXp�<�������U�< ���K�_�\&�{B�ۚ����:�	�lT�ΊQ���`��g�!�����E/f�h7�it�놞�l3_(?�缂.^㝝L"��Ο!"0
s����Y��"����M��,BϠ(y�#u����n�׼c�ϫ����@ţ���$c��E!S1��Wi%#݋�*����+3��e�ŘpNC��wy4퍹�A�94�i�$��FZ6f��ёp����4A� Y�v1/�����a����,A$2!b"(-y��O�h�,)v67#��>Y�E��[�*
�G˔��$�l1w��@�$�?�0m�&����q���W�[p(~N���7�ŏ�Di���MLM�j�^uQ���3%����1�#����*����XTSf�@���9��2�`)�|��*7��K��D��z?�$�ycA��U��^�'�_P�����E������w����0eS�,D�tڹ2�f���
�%o�U�n�R<軫z*\T�_0B�q��p	�]
d���m=�EE��]^�?'¼��}�p������jL$XM�i��i1���
rC���yF;���-�s�nC��-�8�{0J,1��lb��H�V�k�?�%�{	xP��H����������A��3���+�!�L~k�(��*Ϭb�I�x^=�O�t�4��V���.���!/�w����{"7shZ�z�~�j����8�G��Gj�7B��mRVz�R�*�ӸW=	��'F���{:�T�.�`d��ts�0��d��z-��H�}�7�gPL����Ր�l��񮨯Y$���#�?�j�i�Z�N4�w��Ydx`j�F���'2"�w�K	}�d̃{U�>�چ�\���~s��gŨsy"��QYn+�]L��?����:����(V�y^!1�V��N��n�M�F�����������te���B�9�o����L�����6Fׇf�����4,�{��s�^�W��%��BD�)�/%g��4D*�!��@
TD��s�p5wќ�G���7��YSϭ����K�([���׾4�~������"������kַ�Xj�����V���e�޳!֯y #��|��[����s���4bG)��4����u�8�m�kh��
���S�P�(/�����M���!��Y����?�Ovd��Wj����(�k���i[�J�Z��eR/{\D�e�(�f�U�/A�st� ��J4鍆����M%.�! l�9�<��U9Av+M�d!}��M�[�Av�(%�����+.=%�p�M�2��Z%K�J�P�!pUԅ̵�[�K�e��p69��������v���P���5�.y��l��0x��ț�!��6�60��#F�ϙJ�@�8�@{�Ée�悘ˆ�4ܶ|���(z�f��NvO	-�ӟ=�H�i8ѷ���;��y:9�� ���5���K^������iS���g�K�Iވ?�;����3�TR�=x�5�R:T{[Q^�g�!�@������x���˄Nv�}"|���/�˜�P�hU,��[БG�؆JW�:7ų����d"��7y�������^U�#�34��~:v'v=z3�V.����We̱3�q$��pʬ,���i�+J�1��]��պ�O�J|N&��������PZ|4�@[���<������pN�+4������
׏�#+��Fy,j[u�._��3|������,�hb$R�2��O�Q:���C?�
#�!���=�Z^U��s
���G��������3�KN$o��)�Gو������'&a���NV�j֓&�Dl������K�r+u*�����+ư"&`iJ�a��H�)>δ	H�(��eX�[?L&�M���t���@c�{��!�`�C{�A��c^H)�Ź����u�vvsb��l$�H����ђA�0�,�c�>/F���I@��/��$���ԳM	r���f���J�z�y*�O^�v3����C�?����r@Ɠg�@�b� �x�?"��K� �Ւ����|��A���Y'ъb��KS�?R9ٛ@}̨�?4i�p|ޏ5�:4�'(��L����t��j�x��C�a��_�wn���+�<C����z�ڋ���6C��9��,��,2@V+B��KQ��8���Z�؅m���6�R�:ԁ{V�_�v���*�i��j�������ȅ��Q�?��#ڝ)�"^m�5�w\�j2����ra���L��m ��a`\�C��|Ct��Tu�էN/�|*M�� ep:�Ȣ��[`����7��~K(��e���]w���84�8�N��b5�0�J�>1T����g4�,��UYv�E41X��Q�3���cxC��zRSX�����*�[���M��Q{�#���լ&�#���#\H0�	�k������#���<� ϶�8kn�H0��$fi�0;�I�dZ�B0Ǩ�j� �5�@��~��.2Ӆ|�D0ލ��̶^GGX������ݰ�f�K������z��>�^F#ԋ������Nt�KԽ����oF��MXx��>��<D����-t+ͅ^ĸ�Q��ٹ{,+=����y_U�� ��T� �%d<t�3��c1����t1O��M�^ZH��6��2�4%߄<���s#4�@V_�D@�}|L�+,r��3Q.�|d�P����!�TB���bhLbDL�\���<����N*�[�PBL��+�:z��švQ��?��~xm.��[(�2�b��g~!��`�W#����dY�Q��H�u�&���R<=x��ۤK�1mV��ͤ!-�?{��I��>��7�/5!� �f��M�\r>�I�6�R���3��9�V��� �ch-W8mO�;�����0�Ygʅ̳I��A�q�(}��5��=F]��EY��#a ��*#��(�U��icH۹R����z���	��o�P�6�`HW��JՈ���{\�w?[������6�S��4��'�Af��\��MP ko+
=����.���ڻ4Ù
��D�D�R���r�G3�1I

f�y��쩓#���V%�#3M��Q����y�8e_6Әc�\��s�|�����&="�c��~��
���������T��0+�R�+J��Z8Nh�IԵ����`V�XG>}������*Vg��{b�S��;�\�{e��*�d�ņ/��t~���2Ҁ�����/ź�ZB']QP��77����U�\o����B�Z�R]��	����v�4m���N{ts�VO�u�#V�쑽V��}٢����*mv���;o��J�͊7HSc���K����S�6"�y�ߣo�zXj���gc@�L�|{K!���������p�fp]nTU� X�	hJ���A�#ć�g��q�R�$Eo�Vds���ۋ���'��ǚ?7�Y5���l9G�s_ �'��a�p5�|��p-��VƬ"}����R��Rŷ`_Wǳ�}ɾ�^�F�h=%V���H��/�0A��u4�e#�и���e���a�rE	�ipsH�A
��
��m�U�����(+���d?E������IV��@%9��6�Ey�T�o��il$����;�K�ɤZƮ�.���T�me��	!4�?I%�c�B���3ȯ9��c�dj�ıxE�	����gr�E]\�O���i�����Y��FB���ܦ��T.��I����њ�;�$Z�$0
��>Ttz�?���)ܤط��)�S*�]�מ�{��f����9���(���w�e���I�MX�~����)[��fs�W(�@��,+4�K�_L�913�U��ظ�����u����5���xg�~ἵ_WL���Ih�|jSӮ~pR*�� �L�2ʹϠZsD�Ai�R�:W�v�{�h3�q����	�@�O�����rН�C��U��$��[Ϫ����$.��];_�#��B9��_�h�`ޝ���E���:�bv�㧹�*�6�s�nҌ�K!r���2�1#8�߇lg��2�jQ��6��a���[2X��y�@�U�B#�,V�8�=����Ί=�]*��z�`�)+4w�d/��@�ubj!��D��|�������2��Ds���;a����Z�����C�z�gSM��A����c,r%��^/�z���~��e/�9�xx�V�#�S�o��k~��)�Ϻ̀eR���� ����FOG���'M茁��7m�R�jG�N=^(5���ίp�ȳ+T`��xvN��uA���^I/�$qi��n�P�AJ�\dIX�O�:q;���;H�{E\ۣ����>�._BD���fB�����R����)�w��ª�8fG��V3�H �J��71���F)}�d{!rҼ�{����x���Tڞ��]މ�(zA'6(>Β1�7jp"Ҝ�r���@	T��%��f�/���+Z��{ӧaA��dS�x}�7��(g('��Ǯ�ͩD�[\��WQ�7�u�qS���j�p�R�FI���+@�0[lj�Lˌ��q�������4���v0Fg����.�H�,��ƫo�х��Tod�C���c�Ud�����Ù��U�~��)O���ѯ�	K�H�2��%D��r�0�+�K	�7�˸��b�5�p���/�>�-sz���hv����J���D���so�eQ$�97�{��b�yӖ8w٭���)�Cgrd=�
���j�ZL׳A{���%�\��1h��K��kQ�-7����vA5�g��e��&�A)�h�B؝�\�� �}݄��R��wLq�r�*� �h� ǟgj�RR�����	�J�qU���Vl�;�vӔ�9�)+u�NJ�s҅3V�G�
X����?���>�A�f$�ޓiq2�U�ٟ�J��ec E�;a7�A�C#�.F��%��c �e���W���=�5S[���qb���Zj6��#���~���T�y�{�}g�HlK�v��Ǿa�}��Ǌh��
,�D�n�㆒�p��u�(c>�5���t��A��;.O�
�]�f=I���s�z�$��"��&T! ���V�I�2l�&?���P����"-C�K�S��h�X��}��f\n[h�S?o�M�sر�P �)���<�L�]΀p灾��R/�>�1��ZKV(������B�o�Ϫv����ctI�ykǷ��%Q��rF8yWi�]Е�Fv�F����PP�P_(�˘�Wm��|���u3��W�k��d�-̯f�!3W�C �o������ ���;`{K�6R�AV!aX���`H�|�q^��-`[���7t�&\�X���Jz�6�����s�Qo�Ɩ��]�冷V#qC�ګ6���>�h��]�J��ggIs�Jđh��j���$����M1 +wA_şN�`���M��!�2?�n�� ؠ��� 1�F/�8��7��
����q��|{3Ų
i9�h�w�ⲳ��g��@����:-���XS93J���K��Wa.�m�Q��m~�I���ﯹ�bP��2z1�v�[�c?#S���dR:^��A"O8�����x/F�dO�;�Z��3��c�y:>���bZ��ҩ2�L~T�������;��ꂮ� l*|�	w��>-�c�<�v\�b)�8��z����e�/����a<ăPk�����>-���	�fz痩a�z9���$�n��X�S��,��}B��BhUom]��ܮ`��7`��ҘB9*�O�>�t��z��q!���g1p�4ͥ��/� �7xK���A��)c��%��?�����;��.UT�[��u�Bц�V1�>���4:N4���y�*�6ݿ'J�ͥri��d2�O��zp�YmpG�.S$"��^1��	��q0F��F\5��O�I��`��ֳ:@I{���J<C:IkI�^gd�E븷2tUO��˘��90P��t�It�g�z�V����
�"Κ���T�h�:�$���WV��p��4y�0�|=|�Y>c�F�h�5�'�	�d'l~������f�Zv����j��|�(�z0$z��Q��X��������:���n�����S��q��!s7�;$�"�)�n�řd�C-7f��	����nJZ�\#���,Q����s�,]6�}`�ç{���-3r�W����i�����gkD	�����	�x �����C&����!����~�vL��r?B����j5Q_ԏi���������K�o�.�@)v�J�t��/�l�tM5�C�:óe¬��f��u���"�<��mp$ ����պ��j�-¢�?�L�(7�8$�Pk������.��,�D��+̯!���g0�\��OCp� �K�JS��t �e?���?hO��F},���j��'-iC��Q��׌W���zVޡԸ��ǹ�1Bq�m�ؑ��o:���hs&7��.V��"f�;�&��/h1�����q���ݢ�f���ơ�ey�"ͦ��x�M4�d`cr�)`������_t�1�$ɢ��
���B� 1#���<�I��ׅ�@���o{�;?��~7D��E�4ܢw3�Pt���6w$C��������(��t�����U��+�24Z#L(I�?���k��T6~ZKS?�o�؃��F)��Y��\)\_�[���R��^sU�E�Giϐ�)�E���\~������lY0q���S �!�vzjQ�Iᠠ�&[��PI"�d�C������g��J�K���-��F�=L�U�4d�y����$� �$����Z�Ͳ\�A��MG���/n{m�rW1��;ހ�aRs���J���Ku�;}�3aN8�PO��3�t���&VXj�����R�R<���2!�A9����������j4f�o74�K��T5��vn�l���ԫ�Lۇ��Q�(����g��\��	0oS`�G��\ ��cp��+qC�x���jkR����V=`X�v��a�O.1�g1s²����vN����	b�5�&r�oGڠ;�ﴈ�N}�;z&9��;���h�>���V��-wm�*�3k�\H�f^ޏx˔���@��SN
��������Bv$:�,����%�!γHj�N{1G��9�b_>� @�3"H@��o)Qf�"(J#"%wH��k
r7�.�y��I��FI�u�0�����B�Y���F2f� Xds�g6�j�~�0Lܼj%�6�Ĵ����T��܋#���(��� ���u� ���7ig7�-�m~��^���1�;B��`,{���g�D����N�`��Ή3V੆�U���z_���|��Ħ(mI2�ȟ�P1����L���n����(E�C�S�X;�:������t��hYK��!Xk�	��❀��,Ϝs�i@	:�)�N��ف ќ�l'3d^g-c�^βR!f�NBt�5d2��:�i�-(�=iEGQ~	p��{uK���/h�|�����z=�O���2��@}�Y�y��X�����(J*�;z8��S�"V6��5��b�3�x6�Fc>�eØ�Ce�e�3S����/�Hp��jz>��<9%�L:��PE��&�*��?��e�Ezz3D�,_EX�Ӆ�,d�8��F�;�J���jN�2,'!�N|	
۠�/�ؙ?�V���2���3@���2�5[y��23����sȁP����'�s�^zk�>n��7]<�>#
�)F^_ۦ�g����W���3Ԉt
��y� Wu�|��ܠ�hb�C\Y*E������sC����w�H������Ee=ي~D�d ��2{��_��'�r��V���"�����f-ŠƁz�w t����z����+�T$�!�ys������{j:w��7vT����l�ބ���e�#����ʦ���"�����mycu�U�p��2%ƞ�BR�e�T��n�u
��t1�����=4I<�Xkk�^wf�1m�zX��w׳{&�Ks#�3�J@l@G&�N1�y;�U	���<5��>��'~�>���̆��T�1e��1'J��[���s��bCp���aX���t�Iܹf䈨QЁmYb�ˎi\]?�gO�3��@/2E��5'�L��=�'���O��T�g�}juYk��ә��AJ�A����M@�t� ���ve��JA��0�S����ֹ�R������z<Fd��g(�v]M�vsC�J�b�=>ଌk(N�R �a߃B=��k����:�0�A�`R�F<0�c���9`RbA3����]P�!8۟�������G?H��&��|��U��랃Y���#��՛v�k
�Fd�֣�M�)�L�8��k�k7y���U`ǥ�f�Y��tNy8�����X�v�;(~Z/�H�V�Dn ������AY�_�����Ik#�q/�{�1�#�W�aR�Z��Sy�~Zm��`�jB�������j�|P!��@�3��G'��I7�t�G��nZ�f{�}���wB�J�@�>I6��|s?��dT�eR��܄{��;S��VӪ85t�����v�$v�{x���E?�>���������u�����fL��O�O涂�Qo!����Ni�Tӣj�pJQ�圌F14��LN�����g�*J�#�;���%p�M0N�$7����Ҡ���RC���M��/i����ht\9�H
�����($��_�/b�U����G@�ܿ�aO�`$A'F�U�<��4��)�E^�g
�
N=/��˱�9�`�2�9�5�۪v7*q��V(�)9��$r���"-���r�S^"���$�����y�GCdSZ��d'R��b��\��[�ǜ��)�桬�If"X�@٨��$�fy,M�7��m�T��hгU�E�+���œ���S�}��l&�AZ ���}vܴ}0�i����5�Co�6*=� ��V���3��9i��� ���ꉷR��p�����JLZ_��)?{ �Of�AT�ө"]9�����c6��M'<�d/l $���Ĝ��ʾ���Ie[H�m�)?�<M8N���k�n�˃;����Iђv�E�.rG|{K�e�H�#B3��{3�����y͚�93�w=
lq7�)�Mr6�����-$9�8�qt�8�Z@�r��g����R�=�J�!�qq?��۪��H�?(�'~*|5��֣���|͔Y�fԕ�U=�37v����p��io�^�?O�%27)�O��'<�9k�6���[�N�D��R��d#;��$�qړ���r!�4�k��Y���V?�N��
���9�B����ѽ�7	�MP���T�.��`�8o[�m0\2A�V�V!yM�!z���
L�ѫ�"�z�����X?�`��U��@��p�8�x��wt�����ڧ����bm��[��80Ŋ+��籭�_�f�]���Z���Y]��\��h{͢���<�3����T��	���r�fc����^J�t�ߜX2�d��!��5Ԝzy߶�!��l�s��ѧ9C~�TSr�n��QC�T����ȫ�eL�I��I��(��IeIȈV�����0�]���A5mN� �8�r����a�*����!NI�����Ro�U�o��2��TM��yXoI����<2�'�X�B�`[y"���5�'�V�������T��̇�0D���{-H��*��RI�sv͕��t	��#x����z��	�9��7�c��޹>�A�&�����d3��n�n����2xU��Պ��T��=��P��!佔�Eۂ��3��>��U"��!��~�I�jyhnSx�>����:Z�	'?1b�؈��#S���m3B�����W�v�៥�xb��)���J�|��fH��Ĳ��i�&P4�jhtB��5'��Uc'�j�"\��ң��8 pz�͡L����#᳢+����ʨE��H��#�2�E׭�
xu?D'�֖vW�[r�^�������Ն�)k��),,���W�A��W}��XR���^,tZ�wBB�$��_1B���G���װWХJ�y���1�ݟ4�5�s�S�()oJ�a�y�T�Q��6�,�Ǧ��. ��L�V�����f�K�;z_Ĝ�)�oI=>$��j�7=~>��~*����P��zo*�v݌���B8o�%��LZ��^�����@L�>�$�Ά~�r�/fL��+�t�)��(�f�V�o�]Y�D�_p_���\�^�Mʪ�Dp�]9�=|@�(�|�Z���VU'[{��z��N�{M���J��(�g��f$�>��'�?����&�B�6[�|Ȼ���g~��-�hAr �_�jw=�&xFL@렕�m.��1�_�h��DlQ����w	I�\��S�M���{��;B��@Fٯ�&���F�u5�V����|5���9��q~�S�����U]��I !��>���[7z�ˇ PB����4��C��*��{��������'M����K��Gn.�f�g�K�.�'>�Ҕ1��c'-�PU���� +#��+,G��Q>)�V�������c�J"�(D�X�w��T]�
�!�HUZ9Q��4U�K �M̩C�j����v��(6����?@�TeVm�G�//�����>�C��X�^�D�o�)Ǽ��_�S�Bc��Q:B��W-jΪ�3�"�t�<��o���������,/y5ɯ��X��w��c��8G]Tg؏��0�&~p�� �E��|��(�q?�������p�i�3�K�r{��?dǍ4L\~jN0d�\lM8t$��28��-p�R@�_�����қ���j�:��a�t�u�Ax�n���{/�pXZTN	���X�qX��,�F����5P�T$ѫ�'2�պ��qnY?���,m�h<O��:�"����D��!:���U�}��E�$!=`;�m�;1�~<�F򯊿�Gf��O��PC?sCp��q0T_�;X�Jd�{�yH��zV"�"��Q�(f#��T��9Ռ�!�A>�xϟ9�|.&�`i�)����PGKt܆�;Y����a!�*;H3��JP�U�1���:O��o��z0��W��������%)�h6���T���!����/�c����ݏ;�mƏ�,���?�j��6����ٳ�*�jM�S�<�������!d�h�5���{R�:9O�Hρ���><���g��n���?�D ���H�sv9�Z�����6Sq#�4�r���9�N`�lC�D��9��W둆G~�{m�a���*�H��J�]}X���z.�Q�B��c����~�\�RJ6��A�t�ɚH���e��L巪�:V°��K���t��a�g)q�KPf5�)�{QK7�A�/�DE?b*}j����[�:B#\,��?�-�tp[]w5%L���R�k�:0^R����j����q�X��3_���NRw�z�'Ƭ�|xf��(����D;b!#��="�6��E��>,�u'��4N�֏h� �\J%�����7�<yw4h(ڊ{��<�;�9�eK)"I�m����������#k(�y,��(�X��e7���7���n�,�ډ�м&��i�;z\���$�.���_�(��CK�\�����A���0gOH��t;����`ݒL���c�4�$�ޢ2�TA�a� �`�e'���B��M��&c{�̀���.w�}��<)�9UO0N�%�{�u������E�m�>��zm�v�ԥ�����e��&������;i�YR��cO��X���ayKQRIPhG�,>�
�����_��S��RK fO����XccZ\OÉ��F��_,��Dj�R��ȉhW���]X�Ɖ������U ���`�(��0��a�HP��X�w����@J^���i�yʩ� k�fwЧ"�K���WjM}K55���:y(�י�>�p��ˡ;A���T3�~Ƀ<^k��^���]lL���B")gX����+S����[��Yv���8&�n�̷yg�*�WBִg��A���/��ɂ��K��u�x�>&�s�J-���@��Qv�j(���	�O*�UW�](���9�1%��z�7�� �:?�U /�:_*�Hc���
ZxgK�L$*Xi�zJm�Z?�X�P�k&��;���z;*�Uјx�V
1�7i^[���>c���?��!V�{�"��*Ó����J}5�d�q,��q�h��/Ħ'�望i��M5�2K�1G�������dc?��
o��>���,7�U9��"ću�G 4Ug��4;9K�a���/�4���y�3�V�z""dF4�(r��������C�t_���qw�Л����"�j���yֽ
�������iXL3�9E�L��.VUO'�� �<��[q����C���a�����a����q?ٕtjv�������굈GKv��&,@���)KV3���!�����lxOÛ{}�X�f�R�=?��1l���V�H RLܷHKn7W�u���8|�?ZVNz.�ryv,++�ѫ��V�J\��Ѯݛ�Z�h�ܨ��!�����5_��wy�A4c;�M�d&��������v��� �!5d▎�i�(��[S��;��yI��3]֩�L���v+��s�9b�;8�rSs��M���Ⳏ4��w;QT���YG�=h��K��
��6s>6��*f��ufkK���m�]��
��$��)�I\p9���R��/��h�.��Wq\.o����	�ֳ���_~-�Pk�?�}�C���&j獋��T�����.������.]�?e���HO���}���Q��i�!ì]=�&l���|g�
SO�g�P=[$r~�(��w����������H���2�!n�U�3ǣ�:�/e���.h�t)�m-q�#2���Ie4 	�����ƃl
�.��R٫i�0]Ǽ����9� �5�s�u����>���~��E��e�����y��{�ѕ''�%�����@M1>��p�p�ق����V|���0�� ����f?�0��s�bP��E;��h���_9-������_?�pW� �o/�Z|����>�o��k���\�>�R�f���A�5Wo�t��a�a��a��@��`��l��
��Z�J��`W�� >�I	»�D>�����]��i���������&��OـP:;^��|l�{��s����E�ݜ4��j��"��E���񧉷BL�f�:B,R3��W����zVv>0i�q��~y�\e1���*�P��1k�r�}�J`�H���Hp�r���'�r�w�R���M1of ��d6�	ϊ̈�� �V���I�̤͆T!	����jL�gf#\����>�J���J��?�	H�`�t�T�S�DI�\A�Me�=��4�|��!o�#�
*��'9�>i�����f�qi�-Ǯ9C���|��K���+���d����d����ޤ������{U�����,�J��z�����C�%��4��;dJ��+�#ċ�;/�i��skgx����~�ъ�}.~��Nv�g,�����)b������iX#5��W�%��i�{P�-�?��U�ee�+�����w6$���R���9�y)�DLq�"r�b�3��%���	Xȗ���,�΃�v��r���4�H]T��}|�\�_T|9+����6	/W������9�j����Pq�v�4O�	[B�������9Ӧ�a�\��G��E���aR�3:�st,㪮��DFFt���	v���G�}�P��P ��XoAx�2ձ�g��w'?l^&)!Z�7��']��0�D�8���{B�Й�22frC���q��� ���m+Ѻ�F�o���M�s�L5B+[Y��'�ӳ�@�u�C+��qM7S�`e�Ś�Va�+y��1o�'�����@�� O�PHG�bTS�g�20����:܆&z��b�(L�-jƜ).�ת%n��w�4T�>	1G"�����$!�[�:O�t��54~=?}D�lF�g^HƢW���*x��HS'�ٲ!�*J��ɋh-&��ǒ� �L�J>�5k�^�9���s�6`	�o�˚i��)A"4�>>-�4y;��� ��a�aAݹ�H��$�|���ޯ@�a��R�Y+x��V�����+�����c��7��U7���ލ(1D�'Q��r��B0�����M �a+ِ%�k[���p"��S���u�ytM&�E�J�B�뜶E!5��^�(��"-�O.��~L���(w[���;�Br�Oݾh�<f6��>�c��Irc�������]D�!5J7ї���߾��Zj-y�=> ��ǫEP	�����c�G��t��q?�����,����*�C�L<��c�S/������0��Ɍ�:�R zJ�����^��g�@�-�l+���|G�$ȅ9�N���1��k���>D�*�߇�q�Wq=]��GF�mC��k3��nyơ�l0f�L��聍Je{�7z�i����	��	F���@w��Jq���y�0s�}����Q7��@R{O���Gʈ��	4?F��2N�Ky���.A�^1zB���eo��FG�*������^'<@�,�Ƚ<�y<�䤬�2XO�H�[n�=?�G~�G��$d�qᒊ�yx^<���=�ٵve�}�_�j�6�Rr�����3��2���KP����E��9�'և������q#�ds�i����?7�et�*�ů�ګJ���J��5:��o�M���w��"���2@�@O��ҡ�#�Y��_)���Nܠ��Ɲx��]7�.3���\`����s#% Kr�)A�vVa��]R?#Ύ��i{�%��RT�S~Fa+��[�6�;�Eˍ����'��U2U;�:'z����Fih��jMRH��{�߉bŖ�i[��g<;�Hi�Չ
*�C7�|��n�����M��0i%-��\�ת/�pR��%�i;3~�t�D����[nI4�fV#4� ��sc*��	vR�`/����RwJמ�~͈#���(��w�0]o�����
8��"����GȒ���u�W�́�YĤ-�B(�u�(�#Q��<�7��5��a�׻�ٜG����%���BHA6W{+Z�H�0^A�\!$�-��4rj�?ɾ-�9�z��&%��,�t"ۂfX�D{��Z`���-v$���Н���",sT5�;�{�
K�b�]��~u�}-��X��첨pe!>��Q��Ej��D��Wҵ������/<��8��P�HEB��>|J���7�Z~D��KX��g�-�^�`vqX�B�U��H��t�\�f��B�����4�x�[F;U�2&ȩW�����3DE����~�c�����g5Ș��Q*�z�^��;4��s�OkIH�_��v`��,�.�!1�L��#ٕ��>�cH���V�&N�WC��0��Z�� Y��� ��[�%�	�㕇H u� Y�c.��}<`��[W0�ns��"�Q}I�g��4�s<��w�P��XV���!T�E� �*n��O%U��򕕜zy����\区��
�-sm�a_t�\��b%�>!\��?AHy�[e�@� ����%�Y�U�;���6�{;F��n�=G\�kfk�΅��&4���@�����4�@����祼�4͑����X�-ڐ4�ap{��u�@>a��ۗ����U~4X��G[aq�LR�{XkS'^�H	������D:_����u�7+m�e�P�����/��J��&�a��9r>M�I�T���g����� ӫ��
HzY�GA�Q���\w�繼7���[D����8���Ų䖩���c��,v�λ���~���ҥ�6�.��򭩒�8�,I6�Νc��F=��e��a�%L�b����y�2���tR�j�7� #�4|�k����u�sɊaK�4#�I�*c�4=��w|p�n��H0��.� n�(F����d���gb:���צ/hf]�4���8�uܖf�Z�#S݋�I���7g���P�v�D��ve㩆t�uU��r��. ��L ����v_bz���U �0�Lxύ
��5�`��G!n4�h�k3C�`��7����{��z�Gx�m���:;��*Urq8� G�b�Gr�H0w�G��kq�6��t_�]@��b��~�L;/��^����s�zl��ͥ�����#�n�u0eJTJMd���?Oy�*D,����!@V��{y�����y�vgt[�N�|��6`�y��>����o�s���0n)�t�B^{�d�)�&�{���e��kQ��0��I-��a�T��yє�UW �#����!���h�J�m}Y�����ĴR����S5�̀��L/b��#Yq�͞:��$��0ۿg���E�LƐ�h��Z�W���\ ,�"�<�3޶S�DT�:��4A)��.�4����Y�9o��C$�%���.�������ƥc���q'�)�iL�V��e��^�2���� � ��5��l�T@�y��o�/U��߅H~�����|ӊF5�9��&;���f���-F��~��O�+2q�3��v�/�%k���UH�<-:�x����Mc��h+B3v8e�����x�@���G�I�ؽ����W����qZ/M@����
��h�e�z戽V�nӋ�i��h�)����8c��nہ�3��G�32'�0]v�.��ضi�N�[R��-`�JQD/��1����w��OtE�k�E��5�:�w�Mc�,!���1'�r  ���9�Ƶ�w+Q���oF���A����,IR�#V
Ja�'.�|C�^�_���m �+�ʱ�|j��ӭ0O8�ӠS���?Ό �4_��/T�*���4]~hx6j����
�ܔ6�p��)1-;�1�x �F\Ȫ�;��\���K)�[��3����G,R�ț�E�M�,��XRwr��'@쁎I�y�� ���t�-}i��F�i}]��x<�Hc�`~HK[$�U��G5kR�Q_Q*ˏ zH��*s4,4��m��UR�*��+�"��fŭ=D>�!�t�*�9�T��D�No0A6''Q��l|����Z�r��,�Ʉӧq8��\��l�x����		�Z
�F��f�(\�FY6���y=uE���r�\�`8$�źylᗳ��t��'O,m�Hȏ
ԓ�<��j���T�G��WH��
Y���𹺰� ��ʊE��'��=����RD�n��â*特5�*;,���ՙ6A�u�Ԭ�-�����)��W�v��{++���Y��w�~`)�y6J�Ԇ��+`ҳ֯e���1��j���(�f�f���1q��ļ�_Ω�y@H �����%t��f-���t�).vs���(fG������P�0����_���	s�|��
$Fm:ޖC��v B6��"z�TѶ�����*th6À6m�c	��z�X��x��<c�z��,;n�hX�$���5����K��U��
UBEq����2�D��S���*^�wF��T"��7�IZfl�.�&�hg'0�d�t:�`&=�
D���H4Y}�8�	��؄��ÀԦt�]~`����(#dA7��|����fa�or����4����䦭?���t�#�/m<՞�"�4�"��'�uc����_'W�1_�g��.�<���'?��7U#�H"�uv�I~�_#΁��P��d���H�S�G.�\�Y����3�9��)�"D�j[ 8\YaOpb��� ���ƴo<�RT:f���ה�.��VK{'���}*aA�����6R	cp+~���`~��t�ǜ�6Sy�=�l�QV��0�2���G|Smr����ˬ�0���"��j�~;�:�#����e�,�Ͻ�ˑ��e��FʣH�Mh�v�ߣ�����g�4҇��Oy�~���2Mz��.�J������z����Qq��y���E��m�V���o�F���)���ӵ!�W�qt�J�,�+�w�X�EOT��u�\z�L�Apu�;j2��I`�vP
�#��:q���޶,����$ù��q٩6�TGS���na�+յ-
��ԍ����E�Ǳ���~箷l$��� 2r�����B�w
V���Xi�ɹڑ�d���q�Ov�x�]C�� ����yՇ���h	�y����X�[r�߀�C�a�4"��U�s4`)��?�!!�Nг��:?�<^u: �����	7�-Ja$���D��*��� А{W��C\�O�T�����{���� ����}��u7�Gd��l�� <�U7�?'��SPߒ�H�(����t���x(��m3s��Y5���Mx\�C��bv��ڸ���|aNA�l���y��ޗ����G�"�:CFj-��γA�V���=�9�Cd0ޮ��:M�ي��|��b�59���OG\Nt�DA
���"c<ZǢ�!\�d�'��r�R���@�y��$��xq��?�o��/;ٽG�H�/��N�ï�u=kmM�y<o:�9Rx���I��]Vh��|�u!�!��H$�#T�#?!۞�da��u����� /�}{R,-<��z?���:>鴙B<�K�h:4Ҏ���x�֑ޣYv�����$�j]���*8����p)�p��^���MӠ�NuQ*�8�At�M��.0O^���� ��O�_��{4�'�����`�c�
(��ة�8�I�I��-[vrN1�ǔE\J<�~0t߳�8ͅϣ TC�ʁ��A��3 #�s�,�? 9sǌ��h��%j��N�ٴ�l���q��n �Y�#�p��N�WMT=N�H��Q� H�n9��	�mY0�?E��F��e��,P��_��~�{f�s����`;J7
!N��ΐ����&�<�$�6"(	�ǖ-o7g��K���Ѭ0�2�FR0��%���-���f���m¡�����3�hV�.��n���`���:��s�"�6��������~3<�Ϛ[Yw��Եvz�׌��j��3�NWXTO��Ee7��fgw�"�T>r�Q0�o�6�qrf�jB����$ɘ�ҙ��b=.I6�ր�a  ��f=�bg�����BdrU��N�>��G�w�̚cn߱�	���zs�J�vf��B����-7�a�{E��܅'�i�e†�k�����k�hb����u�Q�Od�V����9����e�.��c���J;t9�	��NK�g*�Ӕ���B�bEs�M^�8k�	�,��b��/�f�j�"��*3�B*�0�nu8��EQ(k{��S��{-�������ŭ����
I��nʛ�ij��_G�1�<>��x���5�*��v���'��@j!�ƃ
�%�I:!� yW���j�Y՞��s�dyk���8���0���_�$W#�ٍ�N�,v��qq?�Ł؅�6�n0M3�쐳�\a�Q�s�^�)
z6�y�8���I@���:�3K�ۡh)2ju{�M���D'Pr��&��Q��a��7��QYG��r*�A�srp����wj԰/��ƥ�|Ԣx�3��_y'��/H)�c���5��.L�H�{�׃��ަ�^��.�"�XMX/6���k��l1����#\�D������3�M+��S�
+�#�39�f�*��+�x�F�Nk�u���y�t����oZ��q��ez�i��n�gru��d���(?����۹�)�Zwz������W�.[��TB�T(�տ�3�8Z.�p1d��;|2?��W��+�O[vK���5��o ���V��V��i�2����gЈ�QQ�/��Mcԥ�W3�^
��U����Nq(�μ��9��s�+\5�~L=���	L��#�3=0���Cuu`�tOl���i2����ۄ�p�vq�N�8O��%�#��ȿ#�	�|p��  ��0�5�����:��lg���!]'���C� �SxĄO�?�bZ*��Aʔ���_4���6/#t'>z�����H�,7�����j�[������=B�dRjե�I���oyz���j�)-|"�s� �L�е�[��������-R^Q������f� 5}��}n�*!z��7�0���A؏���,���w���#��.˛D%ۿ���Z�m�-Hݥd���D��ܤ:,��{�϶��<D�����yN��B~�����d���/�VS��J�I����@X�R!��������s���<V �h��Z�s���?/�/�z�f��:,��Fm����$�P2��8̔��6W�l��l����ǪB^'~�,���5a�hK��ʹ?���{�;�j����
2,9�_���q�NkX �3������H�8XQŸ�B�E��r�`�^�󂲋w:�ͮ �m ��x��
g�qE��P#rK:�Uk���(M�j�n3�AWs"�PʂQ�o�(d$WOw�S%�k�1KG�5[.-�� �쪳�]?5z�#A>D%N���e�4Q!��e���P�k�|���uߙ11%�Q���NLX��_,�C����Yu��{���#.[�5�I���o��T���?Ke�ҍ_W�@W),\���,�'#�s�;���-�"տ���P��%�g7]����w=KgJ�H:�G��P:���Z�ώXUvS@ބ��B��V1��MrV�f�����T�T���_]>X��W�x:2��s,c "��R� гZjAXmfx�V���o�Y�Ү�!)-g�l�x!ͱ�ۘ����M�i�?є{����ކ��r9n3��u߆�Y� �:7���<�YI�g��N�
�7n5��Țe������F�߆o�D_9��i.�:%� � ����BӺ ��������d����� �����&���Ɍ��"S[�)��5�����#��S�;#5sk"浗����CE��f9�-a�Ѕ��������F/W`~���9�����V[Lg+�6g�<��;mD��X��ն%�Ϊ���;��P���q~��[t@�)J�i�A�G��ӈΓf��3!<�|OS߆_��R��V��%.5�3�1	�]�̒J�gh����OucJ�{.d�`p��FY)\�~.�}+u�Vr���~�{��x���Jf�4ĸ1��4C9��1�l�.�lO�������D��H%�O��]?C?�zX��
���j¶��P�0}��K���xH�R��(Hu*G�FFpP�`��p�:���7�{e{^H���0�&3s�Rb�Aˊ$����6(�s��bnrK�N߼�h����Q�86v�](!  �Q��CP�0�Xm�'�t�4P��vpSvС*�z�u�$�JS2�ܢ�wy��b�`LdM�H�
&� Ud��>)�W�='�7�H�ʫ.-�W�˥ ��b���[6>0�9�<�5#�[��N������^ Z�b5vb!�VBbH�j9_U�c"��8�li�n(Y#�c��qW>g" �&�S�{��,Y�UDU����������Q^�su����əa� ��_I��}@�'��셋,�[���ヒ��k���=�0|,�zzLGQWs�cb�rvx'\_%�~�y�t�Ŏ�RyҢ2���e��G1.%QSR���%D�B0R��ʀ���m�W�|Bv�j��G��4D�*iG�Sʉw�`6��MFq7���������CaQB]�ay��R���T�ɜ����^|������oF�,�uk��D�O�*��pb�;xׇ��0B쳫���ӣ�[}BT��o�+E[�C�3�*���޼���]d$X�L��w�j��-_=� #�<m����n�wQ��N��`}W(~"�����N:�a��I�稜�<߿T�H��� ��f��X���0�%}թd�,��a��M�������J��3�Z8��џ���������!���������[.1oh�U�C����5�`yE3�j"����~���_��s[Y��q�>/��% ��Q���$1��<�>��U�\��K)�\$�)y(7��^H8�	�bb^�`gF�p�Y��Wb��Ł�z}:a��_tv.��� ��A����zp�8��G�Y9�%��J��M����}��/�4��n�t6�=����VL�R	�́Ĭ6|��X���&�Ha��1�T�]�\�r��|���xl��&��q��f�:.����]� '�BӚ����?a�W�$غ�1sN�)�Y��ƛ$�u1�L���p�{�]�����S�0�܅>	~�ũ�~�4���֘�^��0�n�n�~ځͮ!�������� ���^:��M����`�����Y$�u����֐�L`V�R�k� ��:=�2]��Á��v�a����`�xq��0�&c���sKj,�  `�rѶ��w�6~����D������lj5�$Xb�b���4�J�}�#��x�~��}P�o
�8�L�
|9�A��:�^���^�8��B��$�!��V��h�4��ةM�^�9ݚ������%�9!�c$��qQ�Ӄ�����[W�%���,��#���M=��u��]�FM��\8i�^�_�R�ɼcc���Y�7����$Tc��n$�5=�V�
�b�;<h��3��ڤ�U>n +~�(øϤ/��+�r�x��,��3�(�vU��U�}��p*qx%��5P�cf�4���� �$�0��g�w~e��|��9������/6�⏤�%I��*Z+x6�ZA>|��W;>��T.�ͩ��H�-.-!�0�0Q����砗�32SI�) ]--��@3�
�	����E�y�jW�dJn�����V.�`����zz�S�ա��l����eG��(z�o�m��1af�o?"�_~���s���m|B����Nc���!�4U>
���U|>M�����j�h�q�2h����!!Xv�e�[T2G���	%m�ر��p�?Žr���<z.w�5٘��&�[(�v�L��t����/d���d`��{܌�ԼZ#p��t�x����݅���� F���i��o���@���h0Jr:!�l�U��8D�W�L����*�L��)���v�Т�����#�r�i�y�|l�RXA�}k!=|�>�����C�ck2,�D5yBv|�H�)T���ɛ�eW8R��x��ȹU��Nt�o��Sc��"G���d�8Rɒ]��$3Ĥ�w�Y\Y�Xh��oʎ�p��25:%����y�[�����)z��<����}]
`�������JSz9Za�I��(����(u��Ě��n��G�]p�z\uy�������UT�{c	�?��=<�(��/zvA4��C3�.�>��U�ENj\6	�KG�F�g=&�]�,�\6���]�E�Xb/m��|U	`�5	������l�z����"||-�ݴaX�P��y��4M��m'��S>�p�=ܼ����wo����x���4Y�Py��S߁��Z�P5\�n���_�+�MCl��
X�u���ā��<X*��K�0�	��έ�nG�kq��7�پ<�fι���%a�J8��2��h Żf�ͭB*�k� ���mtFQ��Q�C�5z2ᯫoڥC%E�j$����2�Eّ�t�M�t@�p��T�)Nj$kQ�	>}�r��i\ja��Ƌ�]0����MQ��PU~B
:J�����*!Z���<��_Vi϶@��a�������R�gL?��l�pz��[�$��Ew� 6m�Qw�"��R�ȣ%2x��hB��M�a>�ˎU!'8vܫk�&�m��ެ"TBAx�ӣ#=���3]Nq�]ϬlmaJ[����d	�
D *6Q�yJl�Tl{�M3�A�Û�V�l��fYFR5S���5��P,�A����;�q��\�Ki�-u��� �N�5�㩑�ܙ�2���
�"��"7F;�#�S ����BDǽ�I��7eg/���7b8*٫��^�l�V�	��s~�O�n�B���	�ԋL"{س����z�^�Z�����S$P"��PB�qQ���?�����Ӓfѩ-�I��IѴ�}�^���A��Hs�LL+8�I/�ݔc@��� :��kTK�0�f�z�����x�܇���m-�K6�>#�Yo��Q��mHDL�O��iʎ:)������s�#>@���85���To]o����y�'���m��%����@ƋP�Ϸ�>���}ˊP�S��5�5A ��-H�/�ExLE�ē,瀉�u�{���}�.�`I7B0�V�H���E��og�UI�P+|c#�M�	�=�q���Yi�� �/a�<b���5q,M8�;nйμ�]��Q��s�]x.)�3�6x�l ��N�]��J�	U�8���%��,r-g��7�묎�T�ޔuN��K��/��4����4���TB��y�a�Z7fgί}E��b��V��,�?
��]O�or��P��2l]���R$�#���ǸY��[0K��j=�2�O�D�������V����������\�76��C�9�lC�yD@�L�0'�2��W[E�	2��/2�u���ƣc|>��Ce4��_	ތIz^�,���91�[�D���-�~�rDrZK@g�u�=~o$ =w�b$ׄX��:����k���M�N}E�R���x?��j� n�qK��?�c��YCEQeZ#|Cpi��E��i�;S!��6k#E�\��*���<ʒ��U��i��+J��Y�����R����AU�����H{(�_�L��v>�#~���g�4�	~�g�1�H�s� �Oy����ݙ�'�N����+�(�V�؝�
Q�)��bcG��D'(}�����Y=�C���t���O�a �)�/�
&ޱ�-RNXi|�lvI�j� ��D6���b�iTz�5�Kh� �8�D&h
�6�jY��{��}Q��#s�MI�:�}�ֵ*g�o���Y�����,H^�6��迀P7[�L���`X�UB �Q����S����Lw!}]�z����K�`����!T�\n
q���3�JUB3TR�ϓ�>�K�grI6�:ȉ�ҹ����!���ܟj��Q��Kx�^OݐJ���MNj	ĉDr��J�1s$�8a�4�|ag��.v�������&�#m��w��[����b�mW�Y�e^��,�D\>~%�O���Ɖ:����c�&?;�B��+P
�v��\��	�cém��WxG���P�Qͤ/=v��r���a���%�_��C���B�sQfde��.6�x5�ѝa{�Ru3l	]�&��@���5q����=�+���xڄ�n�]�w%�O�4^1�����5YCr5���#�������JoLWZ�Vp?K��q?���b�ѥ��U!�zB�����U��u�ר}����#�����ꔄ��\��,WM���'�ձ�{��ŔgJ� �f�~�#�4�a�˱���$A�7o��MY@q�%NX�g���(���tY�ͨ�q��eZ��E �Q?��f�����Z�w��m��r;������U4�2�*��Vi�Xf� TD�dL�����@k��F9%�h�Iv7B	ۤ��p�}J���f�=�#ya��0�`^����]Ւh�Zyu�e&�
/Z�&�ۉ�_�����չ��r�o��8i�C��A�T!z5�&o�
����|M �<��QUv���N����S?�K��T4C�*:���U����!�?�����?J�A~����#EY�F���箭��5��d8&��N�~޲�<ľ���B� �&��֦���q��G�G��4eIj=�~e��Д�=f���ú� ���_(�ER��%�9�������"ɬ�W�=���F���v]u~��f��oJjP�f���N�蒇�?����X�%x�%�ǋ{�ѭ8�B
u�d� o�8���v����R��$OP<�eu������l�W�Hք\�7�<[��i'�<��`�t5JWF\�H�P<FY, `��˝�Jt��W�m�잤�5�$M�x���E�ҵ�!���y�aX9��H����P�E�5�5PVB��mu��8���E��ۄ)xA�w|�q&��L8"m����_�?�|���ov�"���0y��E�}�A���ë�8h�N���-��
q�P�%	����D_c�.�l�Pã��瘌ۿc�]�L����e�j�^
�u��"�|v3����P�?�<���.��F42z�*"K���y�����F/7�L$�����ڢ��\������6�
M@S�o�����޶�n�r��h�.Z!�U��d��\?��C�V>��*��ߏ�K��.9�g��B�U��6����z�'��]��	~ҙv�AN�������;���z���~�ЯZ��b���k��6�o�LF����Ln9����l1F���u{�P�#TG�3_W	QD�I?�����
��q�b=���fG*���ڕ�z��#����d��!�����X�B�"��خ1M��2 �'�~
�� >����j���L]��$r�;���bX�OSl����(�P^eE��S�&�=~_I6��&�d�K�@�wf���/½�4���-�#;1���-��q�������
����v�/y�ߙ��~�6��;�=�<�����~�K�v�� �P�<6r(���~Ȣ���(I��|�[��0L�9�I��M(�L��%ڮ���y����~*�EPU��]��";A���)���:%;Pڜ�-�j��Ԩ#a���vۖ|Z��lޫ]�/�Ӧsv�ΤX�ݰ�*Y�~��p�s��a��R���6��)���&��m����5�o���޸�GTQuRva��
gfJ�����O�`��5?A�(S�ޫP�r�	���� �嗐]ʶe���PI!l�v�b�5�����~r��1/���[b�/i�Ͷ�HJ��(�y��L�N|�R$9�B��Xc�R�#��AV����sn�V�@�ۍL��}�<	�I���ߣXo{[�@�,k9|O���|�9Z9��S��b�5��σHe||��=�*� ��?H�k�ٮ�v�tT�\h��v&3:ua��~�yX�W�;=�}��$�Za.pO�S�Z�ax��ۅP��������y;��?nE2N?D"�� �GY6�����I��o�U&��
�^Kh\u�/y�GM0q(�I��aT��f��g<��=EE�Ri�Ǟ�2wq-��h\���A��y�	���V�h�"���/��*vTk!��Eg��͎�UAt�,bK�Di���Ym�k:���b��	W�L�<!hL�%���9ۛW��-۸�7����u�r7��?Xy��`��1�U>�넪p�@J�p�9 ����Fnj�+�0y>ų�ib&K,�kd�C������^ �����$V@���z^W�yiؑ	D6:������@���wzN-�;숖��C���`�\Ӌ���t��Tb��Q�7�N?�9��f:��\�}~�r�=�%�e�$�45 
[=T񹛵3Ũ;6��B�k[�Id�<�ѓ�=���c�MlSh9��k�?qX�Jt5\��E��v���������N2��n,p�i�	+ї	G�σx;�d*ۉ�.-N]�#�I�rҪ�)����_x�f��A�띕I���j�Qh�|����"y�eu����vb�猹�r�哜�?l��؋Mi�o�����F.�(%��ѐx���c��������Z�y��d�(B?'л����,�& ��K���ٛ!OHY��	�+
.��	�B�L��l��p�K�e��b��ϳ�܁�p���^�.<\J�4��"���:�#��E	��H����tgw��%�Kz�Cg�����kDRn*}�F
@��� �a�֒���l�Ӻ"F�������I��)�x�6݊7���'���r���D�"mt�$�nT0d8#� m�XD�� k���)2n�=��a�L
O��!̒5^�(^�R��٘�Ro�Aܭ6��d����\h�.�y�@�"�Z,{$o`*>`����4������LYb}��`"a��ega���e��f�
��Bq��W���[� �pĐ����ز�0f>Y�p��!�@{��7��ԩ=�C�SUg_�ǆ�.`7�
���:S	=�K�M�g�����<"��/�c~O��ҙX�?/r�^��)Ja����L}�qeR��/��'+�f�e��T7��6��Zh�4���'+�2� �H)=�-�FW+��Zu�ݴ8Ō�놰�����`%b渋=��r%�e���P61���Nbzl�6u�PWad��Y�&z���D1��!h�����y���a'.?��4��D' ��3J��K�^־���|X��
����
���c* n��e��oW[�-�S�l �CO7A/�20����o�$�:�kpڵ�r�-ᠺ�ר��qóɑ�4[��V��G�
o
�ʺ o�QQ���y9�ܡ�o0(�~<�ݵ�O!z��$���]���7&JOy~���KBa�_�dԜ��?`>����$Ԧ����Ev�ig~�4��b��2o�Y�a�G󝟉zUj�6s�t�� ��`	G�����^x<g[���\wnEYS��RP��,�SD�V�VC�.u\��Z�FY� ��� �岋e�AX��XeN����۬{2��{z:��;�6.������n�l�h\<�u|��^͡l�yf�n/���5$~h��rƅ��e~���g�ɏ��iy���T�����xB�LK��T�7s�ZA�H�ė-�1}��(w�,�Q��л�����vA�n�p+����q�vm��5��Z���L?b��[@�'�L�S��7���
�(��f�pZ�d��+"]����/�����/�q�H?�Bw9�C�W������#�	G��z�����y�w���8�3���2���dQ[�1�P�i"Ɲ�d'ؒ:Q��, 2���n�!v�
w��5�U��룦|ԯ��M%�*-t�NS\���������LJ|8ٷ9�B*o �c5 O�5�VL�`�k��{���/�	���.�.��̰��;�ɚ�m;��e���1��E�e�f�/j��E�d�eU3��L��7������-���!.�x��2댂eT�{��s�sǏy@���� F����|Z�U�`Y�V����̌��@�5���L�����{mÃ�sf/;���~��'6ՃAT����ܲ�W`��0l9rk
P� S���b���
.�}55��	r��O$U:bC�y���u(*���|�:�z$#Ք��
g��6�*ZVz!b�%]6��N�\�I�ɔ�{A��.o���sT��X� ��xR#�PE�ʀ�.~�OH�kRBD�1b��E_Kbr~v�~{QCm�ˇW�V�Ց�����o��8�DaeQ��|�eo0���ey#j��9Y���%��T�3���?E�N�D`B��g4 ��eb>-\vX�xZWMg���@2�.kPC~ wnE���q ��;4`�R�!@�'r13��Ӗ�X�<jA#��Չ�[�m��]�?N�y���Mz����a6�I���w���,r���|݊x�8�QO
���L^��-Fbt�5'ݹ��mA�lD�r/�<Ԣ��IQY�1_��ќ'��u_��=�ju���Uއ�w�TC�	���9NU�{��g�_��o��0����i��P�
ח�;�F�pz�����vYk���|,��b)"���~�]��n�)4�p����\~�=��tN���Q���' HdjQ�u��wԱ��4p�%�H���԰�@�m��A�/�\��/�������b�)�?��
������<����m��Ț=t������9�K�.��
��a����"�nnb��v���协� ϺD�5~n4'�֜E�E��$����w �Gv�+(�����N�lwέ�j�O�Jx��5�bᖵ�<�u^#��	4�C���ͨ��>���ġ�x���wNt|!����e��������X�E(Y�I�[c���H��6���0� ��i�90yì2A7ftC@ˏl���Ҩ��Ր�Fb������'�\�B�n��W��J�otO5M%�nr�&����.mVp`퀒g|�*����~�B��B����Q��`�l`�p��C(��= }qV�Ӳ�wS7/���f�q� �Ώ��`%���8I��PA�]�ܐ昗e�,�N'n��������`;ˑ�}c�>�۩�e����ne�fj ݝn����v�t�u��r٥�~����ʫ���7�v����g~�K�*N��ln͎�W�:'2��Ǚ�CG���z(�NU�xȯ��𪣭Eu�K-�l[U���ט��M��|�K�B���������H��{����j� �r�8�C(�����Tw7����S���w��	ʘ[���r�j9�����wgw�ʊ�؏Ƒ��sƇٔL�ǚ� {������c%v2��ׂ��zyK:����^����Y]�$V����g��n� Oga]Na mBj�:�	.�ߚ�X�۷�n�+�{�	ÃZ��K��\e��o�[+�j�߄�~���q�i���_�����봍��B�f�]J���,��kR�D������ �������ӛ(���?C��J���4_��/�gu���o`̛��!��(�V^3^2�����}4�v�4z���<L�z��s��$�A�h�����gflI���s�|�ƙn��y-|���F�J>��p�����\�l������=��Tst�qms���?-O5+�ʚ)g��
�j��Iv�� 5ҍ�a�o#]��.ZP�FkC���Y��l��t�'�`oD�5IDga,�l1�GM��f˦�[��;*l��/����t]�������3ʹڹR�^��:ܸ�V��B��?�+e�1�]�rf�&��o�����b�!���qjwr+�]�������&D}��	D�&4پ+�d���H"$�NW�P���ei;�|�IwQٷi"JW�4bP�U>*ZV��+�Aג�yryg�, 	}�����o�E�"���x��Z� �p���(�#�Ew�����̚w��1�K2E�>C;�q\Oy�,���\w�f�ǈ�Hk���.F]ѽ��*����T �?v#L�UD�L.&���Ee���	c6�Y��)���#�c��[O_�I���ڊ�uF��(��xP��ݒG�ھ7�������( �<d'J�|��h ��$5�R�����U q�O��Ȋ3�­H�>���J�7�� �H܀F��8iUkq2	�H�?�ՖJo��8`4���s�Y龈?@�@@�>�<��G	*.a"��d��aJoe��n���F����Wk������^��7.�uX�z-R��1�����c$'de4��g���aJ����
�rn�b��63�[�_594^+�LO5?��`"� uH����P�o�l^�����(Æ�܊�������& ��[��C�ٸ��i��UP��&��v����iځ&\j1R``���D�,(�>�����f+���rt&���T����:�6��J���9�R��<�=�V/��iQ�$��,�h�L��W_�eĺL�Nу�Fe�L�#�����E��d/'�`U�_|���J�s[S��,4�x�w�Tu���R�ߟQMņN����������v2q�ǦrĨ�[U,t p�f���W���sé2&4k���_�s��`e������
�i��F�ڈ��z��0(����P��g���1�>/O9w!��a���j\u|�p�����C}�d� yש���w�K.��wE]1-DVDjK���0y��m<L��n��Y�n����V��A�'4!E��f���@��n��,i�8Q��7/�-��I��Q�8>�V
,�k��rlI������������@��_��0�i>V_�2 ̾���3�:��U �M�[y��@��ak�u��5�;��/By�x=�ھ��V^�-4~�-��o�� �k܏mF&!j���v<�k��J���Pp��7��D���$���K*���^���[��ZB��哝ǔS:��9	}��y��<IOe`���M��Aͩ�D��R᫿\$��;���W�W�*��oE$�D��vּă��q�W�1�^����"�{ր~u���v�.)�UH.�������¬d�w���DS� nb^BM|>��|�3~�}��ΚX��Խ����>p��+����%�֠��e��^���\;�=��!�:G�\���Q|4C�}����ݫq:d���+�ߟs�R��o�k�D�K_G�@��!D$�5T��/6�e�&]��s�G͚�����.uUD����b���kQ���7ݠ��U��'�Ҝ^�B	F_`>�ܘK����qe����z��zk��7�_1��;G]��ʣ�ty�L&3v0<�:ł������Mm�AOi���]��-#��qR� �����}1}��H��1uG�̀�^����7���$�����e��4�* ��`���ͩ������p-�6j/_��ws���k�e_d(��Z>����A��%��^�2��l�ڠL�v��w"j�]����4��X��-ޱ�x�����%#֠A?��y.��$A�Fq�jl$%6��z�P4�*C�Bi����!sGZ���5KwS��/�ѹd�hD�>�u�XV�S�׾
�}U�bO��1_�E��p�T��o�cG:�oĂ��#��>!kiR6�ҧ@�B��F��R�e-P�p0Ru��U}�"nn(PK7������u�T	s%��D��
�ݿ�E@X��s0.M����;��f�09F�٣�bB.w�d���.����$?<� L�y��5��X���8�����$�NzʷE�i?�q�㚆�Ut�<�f#y ]z)��Anb���^�ϊ�?B���I��;j껗���HU��9���mnז�aЮ�	/I$w�OK���5�:�唁�u����
u��,IH����oL���E��\�֝� p�~4�(^jp����,�]��e� ��4קAkg.�U�i2�!'����g�ޢү��R!��D��# 9��%9t�cm��@�� �ߜc[��y[f��l"��9uF�J�PG�;���@h�b4X������z%�������,$��KS�W�%��I�f4S�-*�&o�h���i�Z��L��	
�m�J�bJE�p:�bEC�q�@�
_;r˅���!�>+�1�cR��Fv3E�
�)��ym�>n,�{����������c���Rm*`�m��y��=+�->�6���� l����/Ri���_�wu`61�@��!S�f�;sГ��)_9��t�,e�F,����~����_��1\��2'l�l��8���V���{��#���zv��VIE#����o=	�/�����@v��kU�V�~��L��jCa*S�qDA���TI��nk�T�,o���k��o\eQ���r6�j#S`/��/�l�z�F��9J U�1��f�pE�Zc|����2�D�A����,�?�iuD�����[�����{�����B6�ֽ��uH�9.�ֆ�勭�9�+J����޵��Q���دW��%B�!��Ҋ��h65hZe-=Wq���bc'r���M��l��J����[��%#�:�?�N���~*�~�`�����1mŔF��N���t��Ӭ	g+Λӫ���Iz�Xص�p3YV?'j��Tq�my�(���;��S�R �=�ECk"\�X���x�H�9�S��߶���?�F>���g	�	����ˤN��Ż�&��Z����8�^�����)u��n���;�Tݫ�V2��=�����V׈4sU��:�OH��j�'�}b~F��Ψ����$�n��p[�0�Vzl���w���y���W�p�z�}0	H<L�ςzļ�ߺ(/9�^W[#�-���8Ǻ���;��Q���eq���c8P�0?VY;�{"h�C�VV��ͬ�n�D.��̠��m,��X��T�U�����`Ǩ+�b��M��T�Y�����ˉ�g=��&4�.��=Cyu�"~�o
u���@iA]�"RM�����ת��S��� h4�\P���2#[
��Wy�@���>�����T#VI~�M�|5=3��I��e����]b�@�z�0���K����[�������B�nq���?1���
������<2kJ�E�r$��O��b E�V���&α/.�g��$�Ńj)ؽD�*�j�sRyB��tNӢ��y�:��Lo��J����W�2_�~�Ѫ��/@��La��{�59�GM4�,x�Jy���yD�K����WIt��*�t��
]�s}�-��C���j3C��N'F���ߊ7s��5}��cm!�j-⓷X�uat}t�qM5i�fN��&Xl[ 4�� qd@`;`C
��\}�0�+U_�~N)�sv�!����������dA�Nz�#���%��1����Xm�r�
�d�F9�Z����֓4�9��Hs�<��-8]꿂VO<�?�4n̤�Ƃ�g|_��z��	P��ө�wnF�{���[߁X�?8��d J�=7����#��\d��,���XZ�����^p�;�����	k�
�(��|28GF��ˮ;V��k�U�.q�1;��$=ZF�m���{;��b�.��)G�	nX�+. ����?H���_6f^��=зF�jGq!�e�D
|�N�qÈ?��;[���nfs6�j��~�ਈN��$���r�D�ة���}��?&܄�::�N���lba��y�j,��
��f�Dо�f[��>�9��u�b ϖ,�R����N)�QpZ�I%PA�$p��FR����H�p�7̧�}�OF���moy	�' ɴ����m�$u�=I��2�ـ"D�[Iپ���*"�Ϯ�� ��ά¸6|τ��1y�_z��M�v�}�&_[$M'���	�����	�D�[�؝��N��]z.Yr�e���%��E��J�a��*"�������^�"��v9)Vx����
U�R�O�����leT���o.�t����n"U�g&ɷb{Z����+lq��MA�?�;]��~��-�ʾ��9��q{�P7BQ�������Y�E���v��r[:ry�6���B�JPڜi��w>�'�`�(��� m�_Zkb����-�x�v�h���>&$�����s�Pئm!l*j�F~?�(��!"�u
��zH�������d\�S+�$�ŁU�^#a��0�\������0�dq��Y�5�(�)�Õ�m���77����V{k��S�~Ku��9ed��A��Bk'�j7�TO���vvr4�|��7�鷨�h�-n@]�ŉ;
{�+��m/�(��8�L�v�)������P��S%�UFG�ʆ��6����Ī��ү�AS��:܈�PP�̫�����gPl�:�0��#��6Y8�g�����)1��d�`���c���ICT�_�W)8I�����Y�,L���U[58B�Y�CG%�a��b#���~w�S]�[t�L?�*+w��W�.~�� {�[%*�3M����F�����,�9����Bx�x� ��ёz$.���(i������C9sF�P^|;�T�"���K��kƇe����S��+-FS�ڝAy���5 �#���!���V�h��UV�$��g�9O���օ��9�m��s�;7 IIka]�Sܒ,�����9��IR]Ԧ�Z˟��"��9BP�$6i�c�vs�V~�k�'A��wPK�E��ր:��o�K�}QV� ��9�n���F�1����Q�Qb���@���2�=�L2��X�*v��j�O#�X6	��6jy�݀D����1ȑ[�Z�?!O�)D�FL3H�
�VH�-q�,r>=�.RiS� �+Y��ʱ��$�[�N��)�ئ��t���O����xty�X����VS%z��~��mBE��)�HWIZ�V��+����sxM�p�Yg�xQi�ݲ_Y�;��H:�a2C&zD�{�����C�I��MY�u.(����W;�z����9��GA�^|H�gP���5�|�+j6ůrܮVӽ
5ăcH4�%Z�s���.\cOb/C~*��\:�a�뮥'y7�s�i���.iϕ{6G��w��ٖ\b��v�u�A5�>9�V�SG���ZlM���,fls�JXޛ��6>	������8�S���Oj���_qZt�$���y�6UV+\�F���k�-Ӡ7RY�b���OwB��6�3�x�`V|�*nl�y�] wc�W�p�к��5�F��%+K�ۺ�	�u���{�����G��d9p
rC�1���N�௥O��?�y�	���D0@��a.l"�ugc�u�����ī���P��w�������Z��KAx����"�	=9������!�$���'��aOL�R��
N���`m�ѵަ��jϯ �G��+�
b�"hDґPh4|{�@��(�:#Ƨ���औ�3�W�ɣ�2���J��O MJh�7k�L
�'oky��
��-ZII�C����|�_��^,��b<8H�A)���;�o�-{����q���"�k��*ꃂ���k��$��0a�\k�� ��d7����R�������ߔ�.Q�K<�w0�������`I8}ѕKœ�t��1��o9�Af�����z�)��V�03cX�SЎy��n�լ�T��|�*�����p#�@�j�XI<�|W�EyK��	E��?��Cr��NLH�J��@��Յnsxw�X�݊��,��k���qW�fC�J�܎�l�W�%���,c��`��M��%��T�8���)P{�*h\i��\i�lm�!b�5��It~}x͠��H1���< �÷�S-xW���j�/��Stm*JOW��S�#���o#w"Q���aG����ܽ
<k�$�<�Z�Ķ;�U�މ��i�yH˜�n��.���F�H����G�A����ok:zд�$bo�;��ZM˳�J�ᙉ���5�9/���oe̽!��	��5�@/�ov(���>�$�+!o�N�+2s:��Aw$�e����oj�o	�/`7(Is���V��K�Χ����Ǘ�����7��*�؈���,�[�5˼�x(���	v�����d�0X �D��`�[�n9,�8�� J�k�u��v%���ls��kX�����B�̤�D�V?ʷ�*��&�-ˮ�0+��8M���{�E�J�a�:��C+!UU7�Hb~,Rf��eh���-��n���(��Nl�2�'ܭ���1}�c�D	�[��p開� .?�xcm��Ló����w_�����맇��!����r�_�	��h5��B�W�� ��ȍ)�â�K�*݋y�CbuuI�E�S���s�:�K���� ӂ�sm�����%&>J�~�Qt���粻���i�;�<MG�,J�V�ł�M�˧��k@�5�� A��L�����mg*ck����oem=��J��W���H2�Z>�:���'-Ϙ��?r��#��
��D�a���ҍ._{��a�zƲh�tᡓ��(N�a����M�vN���E��.RlJ�;\������q���+�0Q�I�Kb8�2m����dEZ�����?��A�ꎧC�gk7one�1�"CL�J������RIVkl���p6�Y+�%���co���n��c�g�tz�9�g	���F��v��|�gùh�o��A�Vm<X�/ �m�J� i�D��z���$2��W��d������^���0�f־I ����.�	&yQ���:��޵��d������^ ��p�i߆���Jg�%z���M�񄿏����	wze&ځ��n��]�_��|���I�eD{�S����ssظ��G�>	��:3�[���Ԑ��G��\<�h��⥢�&.�����c�����y��1��� �W�����g|r�q�GL��J$B�DBz�+���v��ˉ}+g�gp��T��ݛc�K��y�U	[� ����pxif�'�- �k�e���k4�e��@��(,�o�YjԚ�s�BNT.d��T�A���ؕ2&�����cO�If1��r��R�ZM�|n����T�e��aF�B�X��K����y#�ǫR?�9A���K5}I�_uty��X���%|��-�!$��L�:L��Ǆ�mϸz�Z����\X��K&Į^0	b����)�MJ9iu6�i�)�>�2�Y~v f�pQ�}�D�{���/�,��\�*`�I�d�Dj��m���;!}��?)i������H9]`V��Dьunz{M���Y6՞�<;�1��8�/'��'�I�H2ѥGbMI�;>!���[~@��/-ЍE$t�tˆ��,��ipQ%�ƺ��H�őn� �X9b��Pb9P)|݉
*��/�A��_:����b"�Gºc�� Z���L��b���V����ŀ�4B�Rf������\�24�gG��!Dz-S��9mT��4���Y%f�;g)�|u+A�٠jKo��(7��G��)�������
K�.	l������)C^L���)֪��nD��]{y�]���.�%���^����W�bS�yk\�~�a0 4�N)9��(Lo`���wy���l	k0%��iq9KD4�`"r��Ё�,�1��^��WZ
z��?�:�̅9�K3v�]�M���6) �ܹ�h.�[@�SO���5B���8��&V٢�F�Y��o�ɢ����R⤄���[0�ڠ��*��쫉]wE��_Uϑ�=��W�鞦q8��bw]��q���P�>V�C��,F,�]sf��7����k
k��$u~�8�M���y��nc  �F��g��}x��E�JX��.�V.���-����>ūU�RN8��UrFVS#��Wr��ow5ժ�G��i%_��ig�f k�Ct/Եxh�A������$'u�C ����n�m�)�p�\� �C��AS��O�U�r���h}o��	m�{��<�|��L3{�蛴�W�M�DF�pmP���pgZ4p����U{r���
�$����7���~��8S!�C�鮓$��m�+�U��H�g�I ���w{+���%�̡M������d���D�L|��T�5��U��ee�W '� t�`�<?��캋�	��>����U��d���R�'�nɝ9ĐL�R{|�?��s.��S�),k�1�W�IK:X��7+=�}�AC����v�h���q� ��@ꩳ�_X 2��ش����q�������u8��m,*�Ԡh�Q���������X���:�8߿o��_��T���x¾����$�B����q;��'?��A�l�K5�]�-.7Z���ʅ���,.���@>=�C4 �'i���n�J��TO���.o�9$s���{)�5.�����+F=至Wn��z���,��{�̈́����T�A2kO^_�W�o��-h@�W|:̖S��z�Z�`.��U<3�AәmR߃{f��6�������9��,�S��!|�7��`Q����vv�#���<:���2 ۈr�,��tB���rVz?���F�K��(��K���o�d8���l��:�>��3�@o��:{� ˪�_ߋ�e#�L�:V�S����%���u(�.|���h�+�O�K�؟�i�F �	�!��K��f�rY�J�@�>�\�T����wQ�7���q6O�IX��Tm|�k���#����t~Lȑ�Cg}1	F�%L�z���n�N��ѿ&3�[�$��=��˷�!d�U%_\ujR򌘾��|����f�g���?ɞ%��{
�`����L߄�f�8��à0L���o��d�NI�C���G�,C�޽��n7d�'R��R���W���d���D�\}��Jz�y��eԇ��V�eY��
��`L��Z��Ǳ�}�\���Jjf�?_\C?$Lؗ��v����ɨaf�T���!�uHѷ]�������Y
�-;d���e�jKȖ,{�q�!�&.�;#��5���j��Tb�QG#�q�R��,�<�b�������������겂�IB��[��kwL�=Df��S�vN�gU򮓥qI��Jj'8��PP�7�Q������W��Y�C[+,���wÉ}wKw|��ё�Gŗl�������w�:�iδݗ��֓
f�F��V�r�/PC�!���-��{�����
��@V��lp�'��X���J�\Ǧ(�v�Lď��� ݦ�_����*��מp;��@x:D����j�f����}���aU}��G����ֿ���BGϔ�+�
U?p��x�Ph3�;%jE�85�4�d|���\g�~�ѳx<�X�J�1��S	�� mgO�Jߪ;�`e�г��Ҋ9�*��c[g�֗�=�.�>I
{����q�Q>dj+�6 m�ѿ�@�]�lY�7��]���@ɿok ���ɢ�
�M D�`�ˏ��"@J����6W+ZB�G7"f$�z� �_��o�<�7C-2%-�?S��*�F*�wnM�Z ���2�p�-�^����;��(��˹A����!�[sN�&�Za�=��2��5*}�Ug��.  BؓUM�r���NH)�z����o�,�#xc�l���E׭��FY*�5X9r�G�l�v� ��ݳ��@e������ׅ�����}�,}pJ^��,6����Y����-rۘP+��n�T��ِ�̄~^�Jf]�4j�[D�a����)��t�%��к~!������t�����Ǫ�b�v|��P?��mW��ҷ�0�ܛ�t�I[#F_�g
�TL���AU��'�Xoׂ�7�+�Z�_���qeQ�S��Y���Y�깡G�Dq�fŚ�H�v�aRvg;u����R*p��<�V2�	 ����}!��4<���b14��ˢ���x��O�V$�c�9 ���?!��=�H��$w�m	�JĴ��|�Ro���!SbW�Sh$�-�	=�@�kc�\n�*%����A+�+���6��!j�rZ<��c�
��j�Dķ�s~Ss��uƆ(�jK�S�	=�?�:�U�F�T�V�x
H�x x�������FM���{�N�'g�Ɓ)����9P�Q�>�i�J�jR��Y�|�CRQ�)��������Y<����v[po�d�=��`}X���X�H$:NR�Zݖk�0߆y��l,_�̠�S[9'�&�h<��8�Rw� ��uZ�R-�Y�T���D]��V'�͸�ö��`�&,Si�/�ꀢ'�ai�J\Tt��<��K0�b�U��sa���h�|t�T֋+K�� O�N��o=�����T.�f�=o��i䃌c��C�-��m��u��`}��/y��"B�g�#�,0��[�#\#Y�M)�0^ �؄X
��5����kp�@��5�*����3��rfvd j���l�n�h�cu!���Ԡ΂�:<S�Sf�� �cFh�p�쏗�pui,v������8t���4l�g*:�|M��6�;F��5��pO_��m�d���!@Q>$M��rq<���L�n�%d����WT&R������K�d1��\u3�T��VTI~�J'�����w4��Y��JN�m=N�]ulv��G��Ͽ��G��q�`]�z�$-g�؜<��\'�7���U���掋�����To�R��=�ǯ����7�J�����Jg40���'�9(H0"z�X"	b�Q�c��S�����STj�t�P$���̟�G7K#�hg4w�5֛�X��/�����]�u�l~�q������ol�G��[���9(咲���g���e"B��B�U� d�=��qh�v���d�Xe2��鿺����a�K�����1��_��/�H�]qc?��N~�b�+��[8
MVn�8�X���ѯ~�.�t��\m}E��GA|م:���L��Ϧ��I�u`u&~_�V��R����T�xf����HI`��(�-.`����_ 5/��5�s��� ݲ\�F��64 y"��'�1V���q������� 0�w�D584��G����F� ��c\/��T�e���K/ ��<H뮠�Х%N��G��)g�>���:C�W�w81[��!��(6�E�1!@��L�A��?Y9d���. �o��$K�}YD%��'�XO�U7 �1&��E�Ϊ�W@F�����8��M��C|TA���[�Dd�k\~=��tA��F6邻�Z6�F�0-�M�R�D�?��kY}0J�*�O�C�r�ǈ\�3ZOߤ��U=�ݩ���$�/e)-,@�W:47h:_v1���Q"!��]!Q���ҌFx�칸����XZ,m�ODFU��<Y+��ｾ�u�܆z6���a�ģ��HW�3�u#���:� ��~n�K��/�;�ex  U������QC���-�>rL�/[���X�q����,a�G/I�^��X���{J0�G��?��eKy8wd�^�O`t7k��<:񣯠+а�:��mr��*�r1*ʺx>�zeP�q�.�wΥD`�n��b0_ь�:QE �m0�n-�P5�QNi�h��bv�.�r�9�~����bg<�9�B�<w2�q>�����3U�i6����n�t'K�Ɨ	���G����Q��"�q~������I+#�7�n����WEat���c,0���p��JkS����+��a�k4��Dyw��a��0�'�M1Ij"��\5���V�Jd`�bea�Ė�ٯ{������ɦ8�aFo�2,u
I���HOr�ʠ�K{C�g���LCJ+'`ͳp�(�ǧ���C�}�����Ƣ�k	��ҷ�2M�l���8w�p���H�p��W��a�A��IMV���Q��#M}`Y��
I�Y�5�=��5Qwb��uc�}5q ���+k�g��A���qF�� ����AY}9�|�"�?��Eߙ��X�$��> ����{����ɕ;�ѐTUfʒV�&U�����ꁧ"��dz�;��������7?�:��e8o��lx�L,�R�.�C�W ��06����jΐ�R���Z;���G����*�KZ"��{���5{RVZ��M�#~�=�Fgy^m�=tly��=���9c���͛��?�������OS�V��:�_G"��w�����+l�=ƙ(�&Ğ�!�憔�e�F�.gE��S�@��mw�Q�$�y���;g�ZDUr��B�q��kk�4m+��Ò�c�g�.�_�[c$Ȭ�g $� �J�����دXau)o����uIR��6�B���.Oz����ɺ��V�����|0����_ON�h#։J
����01Z%���H���=���~�E���Z`5D�^"�nzsC����4���gG���53wt�V��3T&�qB�C�����_�/X����M�)}�.�?
N8�¬�g�A�j���>47��4�g�͈��#�$��Yo�칱��j����5��}�ptO|5U�%L���ZU
��4$����N	P��w` ��"8P���w��;E��u���[p��g��dJHd;��M���H���i�����\��(X97ۮ~τD����5�;�ҁ �g�8k�ZEV���P�07i�p`s���5��oE�+6�F��F��-2f,�S�_��׶b�>y����y��C/��w�SB-�DZ�f���BS�긪���Ɉ�:�����W�4�7 bn·* ]yGg����q�ZB�,f��أ�A�Aq�	lq/H����~��@#=zZ�.N�I���P�.8h��񩺢�-�(�e����Չ�g�t>`��Y��f.2�B�g���\L���ݫ��M��7ʮӉqC�n[��Z�ֽW��<��n^<t������t�ފ'[Q�^oW�Ї�����)�̕g��
!�6��)�U8��,�� �f��b"���z�� +�+���1�\�c��ļ����J�T�AEOv>��0e��	遪�ՇpM��(����¹
��c1\��~�dW#�����2�t׎|N��Y@��z�@�˸���T��=uZ+�kr5�^z��6����?��w���"����_���Y��/���"���=�1���f;��I�o��˪NV����ﶨ��y��1�Ń�Q��B�~,>�cA&�.G�|R?��;��ZZv(��t@ƻz4^��c���Wk���}s�5Z�\�?=���Ο4X���v��5��*pn�,X^i/�~���3�2*�,�*�����;��Qi�yr��#��;��u D�_�m��D��0�i`��HW@v�5�1�A�ϻ��/����=/�V�:����7MV����Q�g�i�!`��ʤhM9��H�$L�K�0�6�L!¨��@%�݄tҔ��>}��Ҳ;]7�5�~���:��W��Ǒn��XіQ_�$��tE|Cho�ͅ׷�U��!�MJ �޲��%'�C�|�r����P\5���Ь��>���i�c���:���}��Tu(R>N��z/J��h\e$���|�b����	G��"h�:.^��g*�#��V�"tm_R���{��7Kγ��pg��I�H�`
�/d����l�-���N\ܮ^%��Hw�G�&�s3#�Y�ƛ�,s���a)x��vg�E���z5b��f��D]��US���M$��Ae� �Q�Hz��W���Y�4���@q21q�[���7{��{�%�J�_��e�Ĥ7�xO=k-|v���Ywt�{KD�Ƅ�E��j�w{8�>�{���,y���|X&�F^`�7� ��5���EA�D�f��yU{��D��%1��gˏ]t����%�Bϫ̒M9[5($��F8]{�����E,D���n�����ũ��t�A���@(Ox�����uW �	�l��M�����
�l�,غ��0Ԏ{qh���Lq��ݼ�܆H\�a������`e?S�s+ͤ�]����5������K��1�ͬ��$�@��5ň�Z�M�=}���ݭ�����#	/�"�H�L�}��]��:�w1����b�<*o����'�[3�Q�,K�Gʶ��#�$Tɘ�������T{owb]�/L�2�
1�|���L���	iY@�{Pk0��'QԆ[mo|:��:藝�*��~�fϋ!�M�JE&��U�<+�Z	~���P+�Kn&���pHЃv	���K�y�oV��P�ڇ�[
iu�zv}7��X���YfT@TY%s�6�[�O~�5h���}�]�0�v���r�55*�o|bC|�������1
R_\^]��[�/&�v? �|�a�@��� ܴ�����͌�J.,���p��b�	%�5e|p���A?�&|m���ӆ%?����CSc_�>'Z�vh������kj�����K�ȨX�V�O����$�Ⱦ�^x�Q�~��!�z�����p�D����70�+ ���!a����\E$5ش��f�F�d�v{���F>?D0U��&��ɚ����|��cS��?j�e����IU�L5�{��7��C�^�=cYTV�bG13�_��gz.�c��v��A_>��V/�'�.��U�dcĢLI�K���e����S�-��1���b��zb[�ǡft�[�֚�b��-�0��N��!W\�Ub�G@�p��4 H�<�o#~�Ϫ��>�ݷk{nB��/HV��lwGl�5E�M�"Q�I�㞄�泳+���%=bl%���6�?e���%���O�|��C��R'#;�V�ӎ���:NT��&����Q��8�rV���D1X��wFY��kc��-	���س��w"`��"f�c��]���qhk�"8,���;�1]��ކ�0�ȕ�c�_�j���P�s��d�7��#u�x�(=tes�����&���2�����k��_�i�5Ƀ_��%>���V8��}��� |�Z��Bb��[�8�ʺ<��b�d;@���R��	W	�}~睥_b�����JF����Č��Kc"TJ4����ʮ��B��B���F�x��<�uw:��:Q��y�Qx��6)]��1뛃�<Uq\��1�5a�=h�VjE@T	/��XK�z�A�R �
'52��o�U���ʠĤ���޿�+��:R�쀜5�B:B���)���-�W�YЅ����Gg��P
+A�,�}t^���]]��E�Q�ٖ��&N��r�F����n�
�K���s����~d����\�~��ܱV�������HX���y;�C����eQ���c����s�`�!���\��m�q������ �^\���]���'�w��+��w�	�6o֖����W�,:��a�AM���W&GE�5�ΖP��I�:��{�r��׏5��%��$���C�)B����S1�5���?���V�$��ϑ{�^ 'U3/ӗ��?j!�Og|�l{@>0T{��n�H��,@��I�@<�K��X�{��#CS2!ّR{lq�#�QJ������Fߝ��	T���I>�l0�n9I��:��[>80�p�C����I!q�����C̈́����x���nʬ
���(�(�� #m5�KHY�Aճ�ޞ���ne��c�|v��j�u��)�J�u���ZQ�P��� �p.|=��:93eO��p�%	�;�H�����aݪ��71�[��O�7D��U�fk�#+ґ�ʫO;O�t@/?�2M��a<�QJ�Ew����=g��頌))�p���PS���Y�R ��pWA�ފ�\�J��WA��z���1jc�5�|k_B L��e2�&�����3s������1�j^}i�6=5�ϩ��5�8��d��'�m>�BƱ��+��Ak!7@�ښEZ���1}m��럾J�˺Jt3|*$� w'�Đ�Ɋ,&�]w�z.��BY����64��35N��){b����X���{�\b��{�86 O�+�h�j��b��m�>(�^iw�w�^���V�*IRaC��ض�`ݕ�M{$D�J!dG�El�2��v}O��V�`4kǚ�Azo
]}	��^F��Y�����qT��:׽� �y��N� ⓾��:��F.;_�^��thkkH�
V�Tq��4d)'����N��!��
;q���3TU���<�-P6���m^���-F2��?Ŋ�ݔ�I9PQ���P��g�M0�m�����,��g�xI]?�h���.C�mk��{S�+Q�;M��Ce�º�F'AO��o}�s�+���6�:�Qq4J�)�����Du��2��Y�FYE+��R�cZ��M��1��<���*_a����0�@L��a�+�4��zț�s؆��BbUV����v���:Ke�>�Iro��#���5�M�y�Z݃0������Q�@Z�l�@H<͛E��I�F�м�����I"Q��ߝy��3�A��7�Z��'�xB''���#Qz�����,�QGЭ^��x��@�G!g���o&KC�U����߁x��iӯ�_;48�Ƣ�SMBGp^4��tl������{8�e�Z��	�7��''�G��D���K���Ś�~�����s+��0!#nV��F���XPj��a"�w�o�
�Vo7�z)��>Ï����3���|�����r~W �
��D�T��SV23r�"]x��$5W�}TȖ�)Pv�S�
(�@YJ�7�c��0˃z�+${�l75� ^7��Հ_�{�5P�[���t"F�X��b��P�Qe~�0���7Ԇ6J*�L�����"���J�{[�	�l����H��ۣlf�	$ZQ�-������\��C*�9i���M	�`�T���uL�[Xl����ԶrЪ�d�j��˴��+��Y�Ƶ`TXs1�%Ϝw���"!�G��$��ƕ+��&<���n����v%�}+������&�0��6��4I�����Y�f*��1��޷�(]�+�V�_���Zl�ws�5#�S��Ǘ�}Bmp�� �+�D��E~ESpb<];�9�R=�c�)m�(��uz�OP6�j.�x��+�X6�\�|I@]Y�=�a�/�]>js��?{���M�ƻRl]&��ۼjkz��v�E��$���9��U6 ���+��2�roF N3v��� �)Iګ߹��1��W������Y�������y7S⊼�DNyh����C��hPh��!��Ut�y�̄,K�K\y�)���3�|$�K��]��Ezi�AzZ��	��W2��^�@�:�RGd�w���K����I�+�X	9���+�v:��'��'^��BknN���	h�D�ˢ���o������S��B�����z��C���I��#�Ú�O���)�b쮲1���cj�*a�}�3kz�a�h��mܖ���1\>���̍�:���.����A�3$L3_�N���X��ތ|z��7Xށ���F�����ʱ���Gǹ�!�5`��r���YqoCg�6`l$��)�6.�`Z�����J`�
�,�fsU'O�8��+B!�^2��'�e9*�"a�Lw���.:�J��[`G�qt�uv�+^s��]�	.��K���u�:�T��0R��������ÈK<%E���߁K��U��!yߋ��dZ�<��liOť��,�v�[�4U��f.�Ʈɋ� ���`��L�@��zo&J��ۙA4!(�Y�r�����ɵ��V�Io��I�n��s5�����a�GB���Wq�J� �K�S�v���6+6SCNNG�[����\��Ļ���|p0f^�o��fUo��m 7�b@���ei���Fu��ܛ����y�gV��k�"�F����:lڟ1zB�H�wgtM�}E���i��8�@;/E��+�h1o�9VU�o���_K�q��{���ţ5x"|��x�%���"(�i4�t�{�o�J�T��P�ȓ�sɭ펏�0�p[bS�����Edvrr����4�����%�ɒS���SF��Ʃb��~'��1��}M�O�J���Ft�q�����U#eR�5�O��OL#20_�H���A
�]u��	�3�D)��=�-*��]�'f�x@aVѼ���d�9�F�ę�׀��\����x9t���FlF�r��J�ّ�da��&��"�բ��T���1����"0w�}�Y�2��i�p��S
�h%�n�BG|�`b*�u��/˽�^N���;Ճ;3"B6�dW�rR�S�?p��,�O�p�[�a�P�N���q�CkH�3�H'E-�/]���'��-U~�kn#+ֳ��=t��Gk��b
)����<�|������	�)yg�1�8�f�N �zGZ;���	����i)�UB�S{#�-�C���Aރ�?��GDj�Ԅ/ry=/(���l���ͬWA��NĜ#��8���FHvLރ�=�|�>ۮ��(��ǃ���*��W��t������B�~�K�h0���mj��A�У}���'$���f3�g+���O�]��uK��,���K��~�UI��Ѓ��4f�pz�=�e�+3Is�\r�V�.ؒ�7IU��H/����~�W`�溡Ÿx g!� 8�Jt�;!A�W�����ȭJ4nA}�v6ǚk��+^�=*<e�ҥ�m¡^����}�0���I1�P�'��^�G�m-NHhx�Pm_l���CRkB|�6�^>R3$*�NuMi;~�N!A{�����O�3�e{�^p�}��7�}G8��^��9$�t���l:��rt%<�.^5}���Ny��[)��e*�*f��)2�7�O��rE6���t��q)x\��5 	'�/�̜�xA��]P���k��c�m8��p��G^�QwU��4$�z�:$=�멶�>.(I�� ԩec�Ψ%�K�e0x�0v�Վx��O�4
Q�_�.�4�מ&�JJ6~��kY�o�~�L�j���w5��cC�Q4�B#[����e8!e�����)3�{ٷ'�� ��祈е������h�A���OBMQx�4�puA���b�#�����׻X:I�B>�!.�7Ң���5����킩����_��O���N!�ߤ��'���Q�1�>>q;톺Mޔ���A��}o��\��fL~�
��JW��#�x���I5��F&�@0.��b�_t���֎�<
|w.��@��'���d����~��x�N	�%L���Q�(wƎ$�^X�.����/n" �ACsՒкQ\2WF!����B��b*I�C���}h���%Yf8�¼ ?>*%�&|�٘c�3���ߡǰV�;��c��1e�$Bd�',�m�"Cϓ�頖X.|�����@�2U�Vk���^�$;*�4�8p�<6*#�g�]x�r��\�9��1zA]b�FҨ��eH'��r���*) ��8�;#�o}�ΈkJZ���7�{����s��]��G��jl#H��|��!��+�N@��lay�a�!A�0L ��Ysd{շ�D��`]�X�.�e���`�7Y7i�����e!��F�vkX8�CO��{�v�s��Ӊw/�
4n2��SO�ͣ�̧��P7�Y�)�=9>tJ�IQ�m�g��<7[� 3,����?�]���5܌���pӆ���VxL���ߑ�+�
=��g�p
LR��|��K|�w$͊͆^�+��I��D��k@�Lb�W.��+N/��� �"�4�{Cq�3���Da���P��F�br����d-s�����:f�+��3N؅�d��8��!j�����<Jto�' �9ll|<��]
*y'�Z�]�ϼl���x��_�_d�Q�����sc-bj��$�##��I��Y�碁�e��C�1��הK���~kB-���Zf�@v���8�8��Mc8�i�%v*�(s�'�a`��}čէ=���i����9�������x �,7�	/!I��-c:[!��ݜNy�oF1�tX�H#,����˦�T奡5����(�f�,ܳ�c���{���D��I��Ρ��Ve�'c�Vަ��3�������Ơ袒�n캳%Z�9p����#N����w�� �X�؁�)��e^�J�_'���@.�l�\{�`)�qJ���Z(��3�ґDb�58��zH�|�zy��#<A��_�&9�ŉ2�b�U���UXQ~$ڍ�蔖�RS������0��hV��?:+E3�v�,	����ޕ�dk��C����}�B�X	�2�,���JA����h|l
.>��A��i�޲Π��z�&|���T;�,NO�{a����Mh��!��
k迒�'�[�9�ʑ��
h��b×�=�����S!"��J\�����7�\�	�m�ړ��k�4s%�]$/����t�φ��z�e̸%����J�X�6���^!g��%��!SiV�@eBj��Z�'@M�_�5���M0�:/t�e�`"�}?��������,����)��+�c皵H���U�>)�|��?��sjji�Z�`{c#(P��W���r?��ݰ�#�Tg����j�2l\t��8�{~�Љ8UC ׀7�ft�ǀ?_���@��r����_���6$��(I2�tȰ���6A�7��x�T����ݚY�u90y���Wo�%����~�G��[[�rJG�"0��򏀉f~Н�$K�|o�:���|-���}%U��<矣u�ڌ�08~���;�C�P�^�}q�ܖ���
�8�f=pߴk�T� Ƹ�3e��&+������-i�e�Kz7U����2N�Y�'�2�cB�e�̼�X�X y��~i�~g�d������.�дT�7 �Wͣ�
��~d��0te��S�+f�k��*��\�x|q�wӂ.RqB-����Ʉ�� ��H$X��e�����˗�;�Ti"��S㶱�T��A�2r)������M-��3�F#ڡ5Al|n5�dk��5�p�sF�\���� �b�7�a:�\/���QbY�1�K�k�=0J���poJ����Y�%��\I5��*��У�{iy���_A�6�����h̼�ܕ%��
u�M$H�V�7�堑 �gd�A�׎�RJzj\�G���J�Z�u���;��o��x�3v����t���G�$�)���#�ᣣy�2�!�P����m.���$}��ja�h˺�g��/�c];"'����P�C��S������0o��lS�d��K/��b��,��ن;[j��v̖�o{�*�9�/ʘ��Z�����i��B����'G����to~�M�]NE��S�5_$��cɵ�|�Q�w
�|JHB�������׫\��D�
��p����#)����6�h���p����UX�
<�`����ֺņ7	jKt��@;����B�"g���m1����A��ǆ������M+������}د�v{"�K��o�AH1t��@1Y���~ZƱDi���b�{�
��<���� �A>�衖w��y������ua)[���랤Q����8M�*f`N��3���1�&R����^��6< ۃ��-�F�LBXgY�lj0�3�7���|>��;袉;�-Cl��_����k>�F`w��Ü#k��[��ػ�L�1��Kw#�ǩB�XۣX���n�3!�C���=�y�zs����|���MG'c�ʺ��MW�ħ��S�ϴs#5E�!�Gm���p��!ރ0]⧋��ʘ#�YE���Տ�����7���ҋ� j9j`:Ȼ��ZpՇ<F4��8��2�AFE�zy~\�YM��0���J~ �Qf���Ee�dS��0���dO����1�W������K�(�̀��|��4S�Y�/[�g�y9�Ư�&zu[2��/0z���!C���t@�*�nh3Y���C�����p=�MfL�Y"������=_�e�n�N��F*�=����(�o��r��Tz�[p%�9�Q��:��>��<�s[�˨Ѹ����U�Q7�oaK@��ɔ��7=Xk6��`��0H��ܲ�3R����c(�kB��Q7u^�t�x���"B�Ѭ>�x d�Q�y�e?y^����/|ه�Du�@B�����X\�R�%��������.i�����K *�R�C�ܳ�Q��+8h�B߭Ț����'�Xcx�3q��#h
��v�d���F��з^6
����2�L�Id#�J��9�f�Жpfpg+��g0��ŉ7t���C�ךޞ�\�uХ�-7�v� a@h��+M 8�ak��+OK�������1$W��˵�VȾ�c\��AT �
M����a#t��@�%1�_�k%W�k�F�O-4Eݑ�*��Ҧ#
�bekϥ���	�=.-׍$�*�e� D��bt�AZB�dx�`�"�Ԃ�����ʆ����z_y�_�$��:�FW�mT�	��<��H!��a@�:3r�8+��߉� ��Zc�6��������_����K�?�X9�]��n�⡫&s�8��ޏ���ő )"+��xS$t��9�U&�C<��H�g�K
>{F�� �g�Π��.
�/�{T~⪩�
lE��Z������1π��3"9��á+[Wľ���/�`� (�k.}s�_z$�A��:����q?|%��X,U��j�;�&_0!�J�(����ww��4�Lᖙ��J��x����f%@yR��������U�Ny� e�Ý!�Y-��V!�� �ɿs�����T�O�r��-s�B�;$��S��Y�y�VO9����d9�3%�(�2�Ļ[�c��"4�a���);`X�Ȩ)��u����1�H�&t/��i��	s�Q$ٮ���G,q�����pX�%�;�J�1�Ԕ�R ��sl�8���#�%�+$^�&[�}��Ah(O^x����Y��3ǆC+r�Z��jKrv䝧�~�,n�E���J��%���飼�����#�>ʙ��E��/����.Fm@8T�+~�s�ϱ9SD���?}��<o��&_�B%pn$,,�2E�@��(/R9z��<�f�BѲ>f��0 i�������x@.��"��}�w�@�+[�Ob�t�=��VR���=>& AU29PR��Z*W��g��*C�X�e�M�h�^{�":��l�G?��_�]�5��\�~�E�mdZHU��s+�� �A������S zF�]��L�	f N�$~f�;IfEG��J��S�$�x:��t�5r_��DXruU��#aܻ��zB	��N ?�I��.#;á,?뜾-�Bb%���`�֠�y@`�����v
A"��;�',m2�x������ˎ��I sh�P*p���r�ҵL1L�
n��tE�6�‖���7��^}<D��H@�[����@o�߭j�z@����x�a\l���g@�֒��M�t�����4{QJ�ĳ��Ł����+�{�U� T�A�Xɕ��ns
��q(�h�K�4���߼L�3g	G�q��{-�֭���b��� +��U�n��VR?�0��vt9>�$8�#ѾL�����M�]k��Բ���"B���t�|�KF/:���!طB	P�h����o��[�´U����F��&����
��&��"�ln[W,�;��%b�r�没�nVn���|��-g�rȊ��=��v����]��:.�x;����#�� �<�#�D��2>v$h�/��>�� �`W&h��ʝ�Dr~��(�O�I�ua_��+�_���|�����~��&�j�XIz�+@��˵!�ٖ'{���2K�����I/�&hCe��F�#����P�,Um���&ɚ˚F��̝:|�L:-{Ǽbl/� ƻՌtU0�^��hY����K�Yޔ�r�K���^�����
0Z<]�[��+�8f�,ԅ�Dr>>����� D�a�����l
c�i��%�~"7�Q�8WG��J��-�؛ս��M���W�iƟD�j6�ő�TD84f��ԗ�[0�Y��r���GV�ϟ�m�(0W29{��`L�K� ����g���*���"s �.���m"W��{���X6�f�r��0���#����5�F�G��|��m�I@2g��f����1|.�91�:�2�6��)JlD����µ翴�M��b[�.��e_&�lR_=�uNenNϺȘ
<�P��!L�ݾϣ퇀~��I��Z8�ۓw,�w���y�Py7P��ϔH��ӌkT9H�Z�b�6p�P�P�#9m
q]���aE��9#����|�]𥸋"�x_0Tqf�Z����d�L��G��l�_p
|a��8���;d�a���x���8�?!��ޖ�w;��^n�ND����U�x{���q1'���*����.Zi���`L�YE������+�׵�AgaQ��=�(����2��
d/cL_��p�����9�@8_�"����/n<u���ӭ����%Ng}��g���+k���9�J��[.7g�)��>1�&ɣ��<�p�+��sW��я��"���G˙�s��;�gӲ�6���ig�1��QL���q�=�omV3n��)+�D����M��_�������(Z�ʶc���a���~��#4���N��b�N^�n��:����0���a���E(+�J����Bk��%�tn��J�<��C\H2�]65���_l�c�@�\g���7�����"��6 ���d!_�֠���?����������n�'��]aO��٦�NT)p�a�hW��g�eGs��a���o����S#���k�r�d����;\/�����m)�2��ͦ3�<C�AŰ�}��� �+�#x�Nu�O�;;l�	%�j��^t�D/�%օ����1}�f�ev������݃.�����p~�^(L�*Tn�e��umY��w�{f��VlI}�[��=�Q־�l6{���SW
�Q����ZRJ�L���u�8-|�M@����@�l�9Ţ�y�`]͇��[�0#0��K�A�^|Q.t#C#U��!����uwe��lRK�>KPu��yJ!�NO����Ӻ�\a*��W��хX~��Mx���m�!f?��k:�B1Sp��V�R�3򀹻_�Z�I�pIu�+s�)��І��F������:�(�XqE�VR�w0���b7�E�p�H]*�
n(���{�8���2�\Y�ܗ<� D�|Waږ����Ӫҕ��\N:pjQ�Y�%������7b��W�3�x��V�)ώ�w�iV��#d�����o�Wr��b���1|P�&�	b(�Pb�R�]W1\[�xX�[�hӱ��!}�7[�~ƭ����
sDY@8a��C��-�ʉE(c<`�M��$�o,s�)zd��b�RLw��A�QKZ�蓝�[<@.?z��;iS�[rA?R5��P�}j�ӈk��R�~$��}r-h@D?��$p|.���DY<�P��˒�5\o\A���at�Ev�/��Z��+�rP��V!��1�t�3!�C��xĩ%y�����.�ޘ{���kM��gĄ�дN��%���.>����4��4BL}���������]�(��rz�h�0�bz��Dz@G{��R~.�7a��O�z�y��V�<��g>�k���~��X�0~��*�I��
h�t\&��(��g�is�ڦ���*Y'��89j�+���?��/FW�%rl�rS�w<�°89!rCK!�I�5ŸE�o�#:��,����&z��(k�^l��r!�JF��PN�a�#I*�c^����"p�4�g``Q��/U)+��irˣb��Z����@H�>#-h�]�_9�M���@�-�Ss٣�SnV�(,.`�hm����Q���TSPK��|B�<{��஺(K�F�Zt'R#V9A��W�?d�6��s��0+-h�y�J��]MܵLV%)��3/[*�������S�<���}W4���W ����T�.G�����O1�F��~\��aVA��Q3����e�3; ��  m��D���k +�B��?�T��M�>o��	�K�r^	r��AV͢�=���3?���W������8����l�?Z�d�M���2 &.N\�A_�a�'��STG��jj1��@�����T��6͞%�!A�w���0��M��x̜�����6G�t�:��D�
X������	Rm�|O�/��SX����*��`�<
p�oA�T��zgc%"�Zs#��n}�⥙K�4�������#��NBv�G���j�ź�U�n�ᝅx��Y�\����G��{`ؼ�ϴ�{*��RR�?�/�����'�X�Z��k��{@�
)_k�NBSd�'���9�ƶcxv�7X���ȇQ�}��������"����ܮ��U�ɰ�I��L4i��z�B�
�i��A�Y��БkˑR��C�W�hH؆���g��{o��Lc�W�����,ePƎq��Ǌ]�p�b�Y���;!ۍ��c�Nns�`�4����a�Ң�0�#�������Ӻ��;��%���:�1��_W��K�s�0�N������E�t���f��G�G@^P5��w!<L1�db?��
c�n�ؘ͙�7"6T��g�}�H�~�g���o�A�Md�=(�HX�q�n�s��{k`�n�H�8����B�>Yad��aB~�m"�H_[�N��R�Y��LD�	�=n$��@���W���
.�՞5<f���;H"R]����N�1����#͖�"$jF"�N�M]�Hs@�Ϊ�h����A��E���� �~��:�g|�-����C���K| �Ģi�;������8��U~S�]�#�Z�V�ij������ם��N��z�.d�Y��ƅ��v�1zq��94��+Pem}��PV�Mw��﶑�"UO7��7o�&���X������˧>ឃե�³��+;�s�R1pe�v�C�������覞"�M�m ��]W�e��oB��?� ��!�2N�V�Bb���?��|b�~�,��ʺB��ݱ��9�
v�3Q���{�Jr+6���"@��:�(���{��*{ak�Ε������@v��aOr�넥���J��X쯸����i�`fL�޿!�\�J�H�Ƹ�h�{�s�=��Du��=j���8�"/�L`;���^h9����Q�F2�~5}v�Z��q��߷�^��t���#]Ó"́�������5t/���E�]e��4ɰ�r�_gg�bt�3��<H��8���ؽ��T����<+�*(E��.�����V|m���Q��t^a��ESΖ��_(梈dt��2�V�����pL�&k�T����[vIS��>8j���w��"���01�9��\76������5�M������I.H2s��q�����T˷���\�Iכ6�g�	��h�-X�w�peG
��٣�"��{l�p=&&�x|Y�$t@��������1JLc�,m�l������J9�8�%
���?��6m�2�m�Q�̿���}��p���#x@[�K/�w��eX��}z�w2�ɐ��C*h��8�>�y�d�f[���M/n
�I���!�z��Ez?�Bv
����vے��qCW�໖R�~�y�y�S��m��ؑo:/�O���gJR)���;ۍsb�7���|�J�Ֆ�@ؿRv�q�E�b,��v��qEk̷���1�nv����SБS��Z��6� x��ϫQ�$��Z�к�M'�⭞�H���o�ua�<K��9�Y�A2r.�(�(�r;g�����xg��D�
d�3�q�S�8����7�R~�!��Lw���y���������A�|�>�('�r����4c�q�rL7	$�G Y>��������-��8�����W�E��-J��mc��X�4Q֦E��܂<Ѝ�dq �ղ��1�^��,�2��Z��~`�G7�S�8c�z��v�Ȫ1�8�$��ylg]/�Y�Q\��:�=J������q݆/���፽���ƆMr��'�g��9 �����?�օL'�+�@~����[�eb�y����$��i��"�$�o\��K�&�6�NN`E<l=D��MI$:��� ��A ��Ǒ��|q�]�Ś��g�ܗJ`�AL�*0"�=��u�f�`�,m�n%�~$:Ã:6+����͙$X�&���XI������m�U)=L:b��}��-��������oH�P=8-1`$2�/N��S^#5
����e�lE�). �n�~*��Ŭ�3�Q�Kw2U�`��	�ő]�b���6��l�ϲ嶱�(�?�AAnu}ؓ�_�ѱ$hQdLj?3ca#���I �#�д+
���Yg���+» 0��u~�w# D���(�Bc�ʅC��q#3�)�H�Έ�"�Y�l-J^F9�t\T����S���qe1�uF�UM�yː]5(i;[:sެ����j?���=�hY�:��/�{��{+7�(�xt�&/i���Ӽ�ţ
Yp�`��B�пnv`�ń�Ժ��"g�:#���F�����Ji���},@Λ�ǹ��^���&٨H�{^�H������/*�i+z�q>;�g�8�},��%0z'�3Q6|P�r�})�.�Z��w��1a����U����^����kT��������"�Ì�&
7s�u����7��Z�si��\8�hdi���Z�(��_ٚ\��)�%-誚�
HA��~�<�ɱ��<�0k"�Y�K�>������tsM�/�2���8�ڛk���ݟ��,5����9V���yH����Wd����7 ;Ngs�ӧ�4�:�
&�Y�f��i����}V-��khXMt�AŴ
K��Wͩd!ZQԗ-��L�4��0��)s/�>ø9F�9E&kN�z�3�R�3�i���a�h3�)q��$Mc>�5c�RJ\`)*V���e�nG�Dxf�|x]�%N6����Qߗ^�����q\��R�◧����<W�GC�*�?��!��4�D�{��t�>l���	�0��yu�v$zԐ?	v���K�)wY�/LU����MBgX���]�(��@�������?��V߆��Č��s��(*0�<еsޓ;�6x�6���?ҿc��(�n�]��}�Я�!HO����$܇�<(1T{��g�7�rGe�Hď�avk�&\ߛ ��kMlg�0�"�X�^R���@G$�x5*�(i������;Ly�)���j7MSR����2�|� s��Cj�I],WM�@f@�&��g�Q�`>��85��Up�ʈ7�Y��&�Xv�š��h��.
�n,�/���}�uc��~1*��nW�n"��NvX��FG�";Yb�d~��Fr�n���B��DB����l�p�pp��b񊂏f�(�r]�K�Q�H{��e��(��8��*�v�8�$�z���5�|��=mN9�zH�K��bv��0tQ����ݍ��vy��������)!y�Z�@�I�q��F����.�J��S\]�&p@����d�(k#�|�7��Ж��	�Yh��]��EV9�fw.V��^ٻ0�^Y!�|�n׋8:V��n*k_+��]4��nZ�]�^��3�K�jQ&���N"�ۯQfG}��f1@�륟I@A��7H�' C7�(����|���,�]���Zu��_�:��������ȑ�=�,�	��FIGM %��%�م	��\�L
C�5.+ң>�#󖔳F��¶�[C8a�1Sj@�?����?.�,p�v
;��	pT�Y~u�C�@����Voc����B�M$����.߶�lD?�tM8���>n�)c���¾5��z|n�!tn�T��d	�K�=&�\����ɨ�Ojo�W$����Jp�5��C�2��Z6x��fz:�S�����f�XF����IT?�|��q�Կʇ�=��r��CS�k
�H����e������Sf��k�0�
������&.m|������;�o,����������Wk�鹫kc�7��=\�W�I������� �=�[�/�%C���R�H��rC���>�q�%'�F�}eŻ�8:.S�EH�� ޱ�a�a ��E�u���4g+-�a�yL���H�,?滣�K7���F����#��8���[�ea�7�D����i�8��2\Y<Ni����&\�ݙ)����zn�'*��,ĿSw/������Yv�[Uq�~�}¡H�W��/���+���,���z4�qW��!�SŨ)/��5��!Z�;{�&�,�.���Y�T����_�x\2,��	�{hQ�Jj��d|�ȁ[3�A��A[6?����\�nP2��Z�%��Y�*��d)��A*8���If��Ty���;����x�$B��4�l4*�닜جLD|o�=��F�2\ş�\�d�G�,�K��-��_A�- eZi�������+�Z+\��D��_�ob/�,B%Y"@9���z&��F�3:3���x��=���f�$�ܕ^&v��^��~��=��U4\�c�c��e�DY�i��nb���׮d��Ia��p�)�;��gZI=}xG	��Ѻ����7��ح�g�Zk����컑��C�Q4���^9�<�}�ׂ���e�b�x��g?J�V���3ًP�
��TNZ9�.�����L �[^����ӏ :�Ki��j�݇��f�����|I�v}>әF{�2��C���G��]8e��DS�E��uXv+M	_k�&�v�^�z���H�7��"1c$�O���3����[��S��7x�'M
g��NB���%i�4E�Ǎ<4����3Ci��K|���#���R��k3����y����m��9%'�F 8���y�;�7���4�e�n����
��VQ�{R)Ng��j?�-W7���QĤ�e�Fv���_�:q��uf-�A΃3oUqH�KU'��I���a�����4!�$�!�s�/�t�.�� 
QLx����:>�*jV^=�������Q�+�L���0��"���o
���9Bf��IP�	��9>ގ=fd�髼1&�{��w����`�_��
�S+N4����,65�t�P~)�",�n��uG�>�Ob����%<о��}�-���ML(4�K��FQ��iRE���5FV|-���7�-�Ϸs���1�D���1��$��M2w"�̱���)s��5!�;�����:��U�ـGP���tBr��9���,33!�λ���W���N6����.+���u��t,�S���ݾ��W xE�9�OP�ޠA�~ݥ��+��Pmڸ��=��i���"�p�E�S��i�D�]Jk���\�nk�P���ǝ %pq���?��x|Bdn��COug�.���F.g���c:��'O���gҒ�!qa�b�%ˍ�v��(�+�L �"�.f����>�#L@�`S�a��k5J�ߞ�]�n�ag�ě���������p_�ԠI��1���W��̔�	&p���K�:�DJ����;��*�D"�ib��5���Ck�l���Pz�Ԣ�temd�����u�[-�OS���O��d�1;};uG�,���ﴷ����/zt��P\����
����i˾e�z�9�^eC����TU�A�ɿ��Y�{�����4%`u9���"��l����S�U3�a�#�A��� D+�;
ƻKEr�A�5i|�
8(m�T�}�
=,˖��.T�MR�E�Nin��.lv��!��/5b���c����P9t\��Q���>h&Ӯ�����[J�w�k������8](�:W���`�m�ZN`�3%���P�5*8���3NIb�}Ƭ3u���=
Z��O��Z9O��y=4�V���8{7ڥ�
�$�$� �����i��'���<Zm��A����hu0����q��#�ª�Y�G�\ڑ�竃�&
��P����LCqW��?�,��
Zto4�q �v.:�W����e^?�P����e�����H�&��AO�M�ǆ������4��}С�`�Yc���gS7�4�p=|�庉��U5�x���wZ�3��$4.Dw6��!�����6�Q�
�"�Ò�a�X0/q�\��e5��Xd7c���q=� ߹S~D��5/$�\�9��ƽ�qI%�q�^ �� �}��<ʿ��f�@!°�p=��}�R��8���H��g��4(B�j\`f-'=���e��Afe
����P��qp:��H�B&��Ƨ�e:gZ�n��<�$J/�E�hU�0�.H���� �Q�GD�F�f�����j�����q�@����Ujd�63��j��eCN ����r됮6��u���O���J�"��y�4{`���`s{M�ɺ�&��:Ӓ��*�]�D&Q�Q����'J�b�Y�#�V����ĩ���!a��X������/��C�/�K'�������{�*������ġG\��jF�;s��)x�X�$m9��������*=�w�[u�� �& �ܲߕ+�.���p�6����MuI��-��n�4�t��,&`W5�ے����
hX�т]��LI��w���zG��g�;9�,<��9�����:&���}�r�ZLOR���	ܱ[Xb$~(�:Ń����J�Lc?���?�s�,��!u����$�hY/LyKj�zR��$�0��������#����9�rζ%� �NF+���_	J��Du[����m?�LN�9�/�5���P��C�$w��;�_^Z�]Gc}�n��g�d�W��4�����-��'������|.�"��J�~��F�JgW�~�"0L��j�ѬZ-��B�Sߩ�7㚟k�I��D���������H��KV�N��Lo�H���2{͆��0q���/�J=����鴎y��0Z�¹��az�Hj�����|�v/ͧG�[�(��.�sA'tb�f����U �Wk���5�[d��7�2Xoj<�-"t�=�Y����(��Px�c�lH�)��B��s8�۬�����%���f��C�*�?������CS�O�l�=K�Ӕ��1�3D�!՞�L�T�7��<��i�̃��O������ɑ�LbP��:�²��O1<�[+�3@q�ɣ�	�����=���H�3b��d��=B�9Wt�³��,E��БyL�k�>���6wU���ڢ+
X�����Q]8Goce`��>e�ik����ߟ`��@c�=g�A����Xl�8u-���]'PS6���҃G�ӂ���<Y>(h�ƊqH�]P���:�$�׭��)�W��<�]�?�e�B�ki5j��4ꌧۡ�X���[k�qM��=������W� ��:^%���,,Z���+"'�E�|v���������o���ClM@X�)^ �W����S���،�Hhc�e	㜳	p!�u�;r���2��*[��L�:�39����~�k�����_A,E�
9�1|��"N�V��S�Ht���J�ur_�1����I��MҪLZ0�_���B���r#�2���.�
�h���3�z͆گߍ	K�
j��������Sxش�V�;��g�5�}�NɐԦ�
����A��b�gi��u�
;7�e��(r�Ul&�.y���^��_<!`_a��Z�L�j0����Rt�f��9�I���B��4�ٹ����d&=7�I���]=��o`�cxE�%�f1���J?��{�RS�ƾ�o�*�&�m�PC�l���������k�I*����N����5rɈ���o�l�Z��={����M���P��xV}�.~y��0�"�.FF��N��I��p����*@�=43���`~x��$h}!A���.�&�`9�,ܡ���o2�֛K��<gN�q�PEB~���[ٸ�7wK���5�k[J�J$����^��H�9��v0}��D<�����K�&�	n�{�xj ��aR�H�a]��� tF����!�lV<��0�@b+eη˃�K�i1�~�\	L�K���ц�&�$o��{���;�DCn��G���I������`a�X���KQ��
�5�FU��fz�UҞH0�<��Y��n�4#V���S�UG�ǿ_�/t09�a�d?6������J[���:{j�����j>Yix�D���%�ѷE���P���9��)9z�7ZV���[w,�H���ڲÌ���[{�����C40]��\�)V-8�?A�)�8	)8�|Xp�e��8�(�^p��њ��O��Ō}����E�����j�8����깔%�s5X[����3�Mϵ�G�Hzbb�)�*mP)�'��l�� �3Y2�y"���9FI�uƬ�;�<Ywr�EA�:�$�j�3�� h��p��-)��n�'8ݱQ�L4��7�4��U��Q�fW3�D��y��,~:S� �,o\ ����R������<t��}�n]=�듽>��m�ƺ����tV}�&����U�C�X��Ys���\{���v�C�P�q���>a�,u�:z��Hva��<a,c\���2E��HƤ,���,��z����g&V�n�$���P��a�"W^��gk��͍�l��yV�4���VI^�ܝ���^��\�vp�:����f�8�FTav��o�ԧ?p�B���	8����$_�-]}��wa�N��^$��:=�ן�2Xd6#����Kr~��eI��˪��"�����Iܓ���I<�NŏF� �e(kJ�/,��i�$�o�k�ȼ�Pvǈ�D^D�t�T%o{�	�j!_W˿�x ��%����P���X�O�3��d/I�^h+@�S�@��%fX�=%���Z���p��3�D��߅钅���jX�ҽd���.6�p��>�����N�rT�a'���t4�h]����D�[���)h�/���3-Ƕ9ʴF�*0|pS%Vtj�TH����7~2�s���|��P�rŀz@��$�������?��P+C}�e�����S-R�޹Y?{��W���	��w��C��b�~j*��Tx*�X~	�%6��q��_�Ѹʪ�Fr�촑�Q**5�Gc�,ui�n�����f�S=��;ha..�1�I�W����S"�h�Z��G���U���D��ӈ,���J�` ���\���rɚ��vy�/�͗641L]�30:ӹڱ����>K-�n�<@@-ޱanK���T<��@Y��iK䍳j<U��"�j��|Ű0��lb5G\��!��	8��~Jr�����?�_�=\x��"}Y$�.�!�>߇�O9h�� ����փ���� �R:#�wA)��H��}�)��[��(z�+W?@ ���_ۖ~9ޗZ<����3r�"5�iV+LcL�g����� � ���ӫ..:�ʈkɤ@�Rʁ�&:��9)A ��Y�[9����r��b�0	�zJ���r;5�Y���j50GC��q���[��g�C&��!���U���t����Y2�E6�(s��x��i�jt�����e�;����u]��}���z��i;���H�����(��'R�CJ��O�Q��b�u�2I.���}|�Ƭb�(YrjC_�O@����<���B��!�U�p
�<-,_v�*|�##�x+�̧�L�ԏK=c�e���Ĩ��`Ĝ%�z(ȷxK��m��a��Vh!�%�h�zA���d;�[O�8��Ak�C�.����e�b��X��m/V-Z�B�nl1�[���!R[�<�cӋ4>��D[�z.���"r',)�t>�֟���	$�<Q��/�z� ��I�Y�p`��to���jN�UˑiR?"e�K�i�Lm�d,Q���.ZV�  �:~��'NZ�7�k��|X����)�f`"YJ���1�a۝��|=�a�;_˻JH��.�����z`y_�u�S���\�S ��zA#���X� e:.�)�XX]�d��REP��0ɇ���`���GͶC��j��h
`E$��a�S��
�%g^&�������b���
YI�߯�PV����+��~�W��ؑ�bT>o=cE��u"��9���(�z'GvRC�e�X�	;JQ���&Υ���K���Cb|Q����d��]�$�C��ި�u�<gO�R�65����j7^��T,��vu:,ә#������m��K�F3���D�q�����^�7b\|������e�0�VL��
rǲ��8zK ȩ�1 �j��D|��6ق.
�v#�{��9o���d�gwo��>���Au*- s�?���k�B���Q�7R$W��M4לW3F�-�����*н֍�9�	h�m~[gÓ��67)G��f�,t`�,�q�b|;�(o1a ��[��� ���M�O�٪,���{�Q.����+6��"�܅��l���R�w~��H�E�|�+h����������a����Yv��5A���,w�m�FLZ�D@�-�?�(I�vD@+��썂Tke���8"�VO��腥��OW�IAQ;/�q��1��:���� �q�3.T��'���qC~/@H��<OFBr1�n2|M���B;�����|�pK��������x'���Wh�Ӌ��dC�S�QAwʀ7����X6�Ϻ�
�1S@`g@U�o���!-��V�:/�x�_��Q�
|����o�UtY�"��8)��A�3.V�i���-"�"J�T�M~����u��(B��;9Y��R���D{H[r��9�jĬzPz�?s��	+�28�3[a�=0S���\��\~���Br����4}�Q�$�G��H��[������M0,h��S���2?3O�x������+=J`d���LmT8w`T��B��L>�r��ĩ�ûQA���Oi��K�m�2�MW��?��l���a?�޻t���(2��uS}0 RN�['kX�����Z��![n��dm�[1���\QU��a�Ӷ�E��P���*�-L1+�~*����CQE�b��)%-��X�'�;[B�\2�ע�@w�љ=r����V�rMe.|0�B�2	'W"J���nk��q�S�%[�"�� �Ot���0�v�x3�m�͊�� *wKDjI�W��0��ҏ7�Z�
�ٿh�� KP��#m�t�L�����@p@jώ0�I�D���bW��2����Ej��'��� �6P�MM[��~�;"�0DJI��?pc��p6�|�7v	�^��(����%��J�F��8��m���A<�ù�'�����N��q�3�;���u��j|�W����|�5�*��������-_Yt��9�G�Qx��[U�)il�x�me%�A�a���3)�<�_¨/�d��C��5���c�n�\��î#��/e-��*�&�]7`��RL�t����F�&�fZ&N��U���Ty��o��^~Q����8�)���l��#&dlMH/~��W�����`D���8j���0vGE��Y"1�,�RA1d��|$��#{mT�)�G@�2~]r*�fi���}R�S�$}C�$���3���k2_����b^j�U4��"�:�$����y����?bM��\�Z%%����,C�.#�L�t��1�l#�޴�^�_���%e
���>��r�=���+�Y�S�A��Y3m���*A�hy�RC �Q�o�;�3vGTO�<EЦ('�Y����������9��g��r
����{�~�	�$���� 5q�t���0�nh��`N�F���{�h�. �Y>X赞��h��"���KPK}ā���"������yA���<��8��w�:��p���2�9g��� �TW�u�[B('�P��r�w�������|ﹰ�k�U}S���o�hԭ���'A\zMf��1U�Ĵ�ˮ�P��*�g��aƼ����+�JZ��U�T������A��C��Y�Fd�4�	�	M.��O�|3������D�	|i��	�$]�D���i�:w&�"�V/4�+'f�?���J�o��(�~�KeFi�Wh_8���_�� J���*��~;4���k��ݦX��J��Hu����Sψ���;'���Ɋ�b�_]��]��$�m1���ڮޯ����>tfky������.�
i>��cH�K�{T7��#��)�BӘ����[���ļHjZm�X��r������W� �J)*Z섺���wFA�b��]�߂�h��B7i�ț��`0�0
1����!�fxD�?�ٖ���~Ip�Ñ�Q�iX��SKJӱuǉ���ޚ8��Q�ԟ=ΘR� �:fX��ds��|�8��X,�ͺ�7%��U*��̵nZ�+B��v���/�gjP�CJڀ?�Rt��z��>����뻱`%~����ƣb�=t�ӉS�Y/���xN�)D;�XAʪj$4T��S�o4��=f���^}�tܢ��ZA-�րUR��ٷv�M��:剋#��ἲ�}�)'RVG����VUK���.>_�#�w=�)�s ��q�wx�9ތ��>����4���=Q��$��j���M:3l�3
���O�H�N�ws��B�N�-������~k�:YY��aSf������hF@])�~Q�2vh�C�8�OH\D�S��X�\&:W�n���~䅁�7�8�T]�!�`2B'���it���2�.r���X�ml6��bl�%�i>��/	f.`�#à�!�^.E��|�T�;�u��d�x`�Z�HV�H�0 �L1PM� �=��򆧒ـ6�P����C�@�7��V�.�k0: ��ц.�\�M0D�_�+����p���u��C}�w؉����%|��ږ��J�-�#J*z)�(u�eDR������F�+�?��
�ǅ��)z�|��n`%��I�f����hS%�I8�C��@�UMs�X�ݓ�2S'�J�D~�A��$��g٢K?����q��B�t���
�4(�z�1k| c����l�>�?�eg?U� R�9�������0<�AC�H6hL�Is`;Y�c�h/8������>���+^��8���m��Q�(a�nD�a�I$۬�m������,��n[��B����@�G�V�B�F�A�����F�{=0P1&�Lŕ5~��JԤ ���ǚCC�"j|Զ�۲y+ȑP5b�{&�ꋋ3�I�]nNg�Yx	p-Q���H^�0�D���^2���'��@��gz���V�2A�K�@���L2�����2j,� ��d�E}t�O�N[������s^\�����'wf�A�e�&��Y�o��-���C�@d�ޯ�vӞ��DR|� ��P�9Ȯd��U���A����q�|�'���8@�c��Q�/��̖��Ť��n�E�W����֨{Ҁ�*�	Yw��|6y���իp8LU���Z+T.�_v����6\��Aр��'>2�x�g��dQ�ՅP&j���d����Zv�,�����Kb��2$|��PK�Ï��s�E.�C�w�h�G`�j�K���,t�ޖ$ucp�e�� �O��1{r`���59CP���,�����[��<Ь�5�0���`�%�96��)y��20�{�qƀ�h�y�i`�(_��y� �S��mU1 �������a� �����J��f�l�*�a��ڷ�XB|ñf:��3�-��[!��o��c��&q�	�$)�D�s����v���_��u�H:�Υ��ObIЧ��.��G�>�ʱ7���|.��'i��|��-��xe��t_��:.������l�h|
Gm��Ce�D׵���[�YA8����
�s{���MJ���(�^�=���MP����%��`&�3��E�et�k>#�`z,;S/���r��O׌�7ADʓ��2�$O�p��m�5g��֚6��I!s�>u��I�dkD	�,�I�cQ�iA8�W	���ؖ�J�a��%!�f3��7��o�er�I/�ܥ�w�"zh���:��{9�\��no��6i	"�h��H����i���P�q�<QRkT���C=�Ok58CAGUg�XN�j� 1Y��O��1����Ƌqhs�b��� ��"��g�$|��Mc�'��*�.)�^	v6٫���^l|�uw*���f�BשE� sP+B�c�[����nl#�� ?��d˥q(�!66�+r�ٟF</J{��U�]�}!���_nN-� ��2�.���Ɲ �<6�q��p �����Je��<��f����fpG#H��4�D���aA��Ůރ.�G;���U;�o�n�YCJA�iP,OIiP�g?�O-��΃�[�țb����S��-C�YoOJ�\i̍�t��@uB&N)}E���j;�M��5���M3x�I"�q5<����X*摰41LSM��ܻpGDP��dr��o����}6��HtvAvِSW���^���rީ]��{�M��x�k6~(?��|�Y�Ro�`xDnM��$�~n!44�
���fC���n�����h�s��X9,�Ԕ**�P�o�_�$��8[<0�=5fL��~�έ�n�I	i4/߯��MF�p���j�F(��bV�%֘dJM�d�����n�!d-�ޖ��d�}K3����V�C� ���3[�ǻ����/�C�(�wXW��§ē��L����n ��y�o�Y'���D�j��Jx�[�SCF���$
�!!��b}�.�p���k$v�^�������m�����4��= ���4-ۄx%򉆲���M��-�'���67JyB]'�_�*��<��%���o��Q�5-�N��`�Я���dBv�B��O/���ٟ�o�q����U�.�F��84������d�����׼>
pz���k�=e�c�>%�M�;�
⁛z��
�оs��5?j���PJH�d�.�&�wz���Q��A�������#�������kHI����}ND�x�B 6��=�h�i� ��q0�&�s�v��>ؒt7��]p�a��?�-�֥w��Y��qs(�0�
f��3�c���I�a�)A�>0�VL�S����z���7�3���k ���3�R�U�݉n�5�Z����rL��=@�ڬ��wr�'iX�6���K�C�z(��F`�C�6�/���đSW�@�觍vg�)�WF�m�5�B�¡��5r���rX?d�ՙ��m��ɫG�̺�{`���v�so��ǃh���c����(����>̼�-���	�j��~ ��5zf��J'	^�����{�WĤ|��fq&&2�@�A-K�X��@k�J��0���ˈ�� ���ڰ��ŋ���4��C�ahU^Pm�w��Y�|����ܸ����6z����/�3�/���9I�^]6ݡ ��ScK�	35��*P�{w� ��	�Nv]�|6g�<-���ʌ5�b~�*�̄^UE�e�Ր˙�G�0㙃���|dg�ވ�4�ʽ��f�v�6����D�L�̸6톹Sј��Q%標w�I�,?E�T GoZ,��?G��&�\A�kY��x�%*zj��%�F}::�|̱�]�tc��5[�an�
�C��m{���m_"V~ϚDs��>*R4�!�S�S[���)��eQ6A�DA&o�����q`�i�e�f�0h���+r�N���suZ�]�B4JUi*N�,d5q�<q�CORr{���N�ӭZ�i�7Zw�A4y��P�ϴٰx�zU�Ʃ�n�1�7�fl=�3��U�(��EO�X����Fv�0��O�'����ݞ0MA�/��/��F,��k~�;������⺱+��������Cq��&���A�+��$�괞^(|w�7�l���xp�xԪ�Ѷtx̗��R[UX:��y]�R<���$���d�b�����tB̭>��"w�����:./�3o=+��~�xo��\P��k�&���$���W������r2�Cg�F��;��C���X(N���=�Ka���� ���I	�ʾ=�`&ä$�V<���4a�M������a7�6�Gխ��[-�R�s�%_U_�<{�����-���J^��������G2k+>�����o=�q�k ��ˣ��C��zX�Y�4B���\ar+dַ�(ө��`ڃ�zV�(��*s��&M�S҂��Q��5��˟k����G��eLq��C�a��@�:� ���驛�=�(�Y��{���=������lt���:>o� f������6D���"��FAf��0oj�SR;���E��e �i�'OYN��n:��x�w/U&�՚��NU�����ه�T
�`^�w� �$6�K�N;���yM �%-�����{�tt��P� ���M��r>xcHV,��sPF��?ZG���O�_����o-V��{����.�`]U�F�pE9A�K�_�-8�~��p<�B�!���b\��'#U;Ӵz��d/d�ɶ=�F�JR��2`��~���?wWv�K�dե\''�����Uɇ��"���tsҢ��z���Y�ֶ�-�{a���jߙ��O��%���.���0�E=֔�u�z,�	k�6 )��r���)�*j����$R�)QcR7RZ*�s��G�SI� $�r�r4q]e�Ĉ��"�7cӭ{��:Ĝ돳<�EYZV{c3��T���]��>�	]�$��_u����W��#Ӌk�f���'Tm�F��{�Z󷯆|�!�q���2
m�P_���̩}�a��K�Zr�6�\�o�n�k��?e�d$C�1�ŦxA��NRs��I��I����ſb�y�������iYq�祾�����J�ڈo��]�{�O��XYs�'/�VIF�]C1f����Ꜧ7s�m |����o��*� 6|�=�ZU|Oz��Χ�N{&(�_M{s{�W��l�u�.�oX��X�a��W�b�����>�#�̛�FVt��J�ʪ5�QZ��{����j��\d�iV~��[a�u�M��3����?��ȗ��9Jx��Ej�܍)Að�أ+�7��������k#˃_�"�&�����9OD��6��v|����� ������˚�k,�z�'Y���,r���~OI.���R����H7��?��6��VR7���[�����9�� a:ɳA�N_a�.v��C����Tz�`���p��]�m-�$=z������n��e��t��<k[#��X7�M#x�쏂�C�Y��̒	�y�d��̙e:�h�@Be�1b�ZC��rXB��$K7��k�,�׳��n���+E��y|� no�ҥ���)�Lt��~}?�e*��r=�(j���Y�`+��;����݅�b�Q,�Sz��9OǇ�T0�q���,]��\f5�ܪE�'$��@��Ћ�!�{��Ş�R�m�'�E����"�����r&j�%����V���|�$�ô��	"���p�/F jܸ��Vn/q����Iش�Z���>��/����q�C��-��rGp�Ft�a�<�r�=�3L(��-��>�%1��e���_����6���kì6�%4����#[ڹ�KY��+��5�;�C?'���@�¿y�ϳϿ�GN	L�l�`:M�e^���%B����()��7zw�zK���q0��8�B����Vh�m�dh�-�3�)a]�[�.l�4�~���o{&�I{A>mX�A��C
8�1��3��D8��B��C�.;�vw/�����u�68"�q����.GI��f�E�,�2txm���<6G�j�}����5���!dd�R����k1�j
��-W�5�S�Ԗ0���TZ]�a�\�< �y��N��2~�d}݋L~/#0+��i�bX��T�HĲ�T@��`r� c�G S�t$�V�m�_��{c�A`v`P���_�(��7l��5��%2�<�^6BT��kVp�]*1�'���.���ǰ�����VZ���@5�$��~xa��s����T�(�0�ޔ��qR����?h!�T=��Ri�7��|��Rˊx:�ԩo�@%�PURh��/emzw�� �t��T��
�k%�����F���,�E[�'� ���$��zδ�ԡ��<Pv�m��.�Ou_�5�Xx���j�q���c1�F����+	��a�w��%�V-��:p���D&�0c3d����ɍK��5��X�S���G^ͼ���E��	��-�NI]Jc�G�J��Mа��R� �'��'���!�)وӢ���/s����6��s����}�#�QO[�;܍����� z,�O�N������V��O.��]cg��.�\��,�s� _�q)Sn7 �/�a�i7}$�z����}��@8��"��b΅�c�4���`aM�'��]��z�}��e&����l$���_yǄTG�ݩ�F.2��"�u��D�7��p���7v���uZ�myo�ب\���,�vHv{���4S:��4\����IY�������zo}Ɵp�.��n���5��2�>�/�/3����ڎ���$Ú#<�2g l�լ_T�@��-WU�82Ķ��*��H��"��͋�:^����L���i=��8V���/N�I`Ə1,T�B-��ZȾ�!e��*��~)xM�T\%�'�ی��:j�,�ő�e���#�Vo<0�c]UJdEJ�e�V/aCI�� ��´%��y�C���W�ߓ,����X�pT�q�ޢ#���lL���}�/�wm�B�e�f-�4��iy\�}iD;�x���V��H`�Ğ��e��-�ÁR�oh���̑q�UQ5-�_(��ҝ��P�3k)�I�tPP�X<���'�ڨo��t�S�p�m3H'�Ǻ��w�G�
o�`[��?C���13��\}%փ����������G*[H���hy✙KӘf.�֭J32�yKs ���4��%���*�N��*@p������t5�� G�KK�eD���I���f���_��s���Kt�Ɠ��`�<QvJ�D�04{����)���^���?�M^�#�g��f�a<3z�b�Z�u�*.�kAD�����и0��;���!s���m��{��rR� �g��z7��4x1���	�T�\!��'B�_��'!���N�������~Jİ�Rct��⻩��8�Om�%�|�K���Tb"�Z�X&;ִÃP��i�8��*�6��i�/��ӋK�]�iH��?<Aq����j�;�"�<//}|�i1�]�}�,|�ҧj_Ξ��s�b��\��,�c6v	��e�X�x#P|b{Q�v-a��IԌ��=��\eZ0�Ą��6,�|Hʳ�S�
����*Y.�s�Դf�'�����߂��RV`��8�ڴ/�dHx������������:&���I����Ƿ��6?�!��YZ"2�ҍC��fB?���p���\�*�����^ڻ H��f�� �4�r�N�fd��iW��F�Ö�!"�EBKU��_��'���C�q�??( =�,�T�� �4��Ǣ�Ӭ���oj���U{��JZn���2x�SJ��{��3B
��bm�bxW��2�
y��Q��ؠj������		-��+��,Tk� "�9���/�.b�;����Sd,�W�S���k,f�V�$ݠs�^_�ҖB@�a#W�Ϡ��u���&tx峺ڌ�
l��
�s$�k)�S������)q��P+��Xa���F����Zn�]C�no=i�T�%w�U��v,��X���}���^���~.�D鸒d7�yzE�x�mQ
�h޵:�ų0R�i9\6RX
6���s]/>Q��wE p�w�\5��t�NU���@����>+��Ng�\D� ��e��"����8'�}����VD_���k�F�}>��C5ڛ�v�|5��4���D��D��Hl��T�'�-i�F�2���{�6��
�]�PR2~��o�o�3ę���V�cx�5�[�[с���//	��`n�2����+�	m!���(p��'�R7!�����`�.���w^jXi�$+�u��=���4�5��:7�6��=�vK-�K/R����{d��EÃ�Я[��C�8+���%�B�s@v�Ɉ`!��&)�A]^1QR#���>�s_��� �ݣ0��<�4J:2)�U���y 
�d!)^Ա��y!.�5�H�i�";�'���('襫o�B�j)�9��<>IĠ�����s]�5f6ؐ!��m���b YLץ�-�X� lpB:2@�xGHb���FE���������W�W�b����;R�'D�',>V�;��{�
�pM,�p��uE4�bƥ���S�� SE�hs�&��$��	�.��up�)���ǺrNH����aJ�r�2��j\��x3�G�Ѵ�A�ΰF�D�PS�,�4Qv�8��F�3'�������sT�z�M� A��<L������{G�^��`O�7
N�_� %�"8+R%�d�/'�\�V&�N��K�o۹n�|�"*#/0��`�`��5���:�w��*|����M�v���	�5=h�2.���N��3��N#�6��	8ࢦ�_��Ifߨ�j.�Sj�S\,QpG�la5�z�Hy��KV���8H2@�d����~������tr��B��`�y!3p�ZTRn?Q��b|�qȉ���h�<���ОB�F���>���c��Aq8��E�D�F.�x߶�Bvfs�z�;n%��Љ�dͿ�/�*�q{Q�/EYxX2�=ڜ9���l�y5ՔH
�:����ef~�3��ز�������#���j�e��\�a�W��z�0{϶�bm;�E!)� ��rc��sA������>�7z3v��N���#�p:l�B�T�[2�u�o�c+MSaA��i˵`�[o�:�ﮝ�����3SѺ��h�c~�!h�~��tauV
�Fd��7-�k0���[~s���.�h�(�,Os4�CZ `���?�r`s.�dk�5�a���S�p�e8�QC�|91A�,b�Ϸ����*hMQ��4�;p���x�*˹I��=e�u�I��cֈ�uaV�ô�ڏ>)��:^��?H��8�F��_�~a��<����sL�⬾�fЙ�Y��%X'�uc��2���^�?���-�#% �[Xڥ��3+�Z����)���͊
6�<���A��ק��Mf�`���� ���xc��ErZm���xŖÈ��N��v���t��_C�J{��N��k
A��ك���@�����7�b�Hp�B��󆩁�Z9�;8<�~x�g����{���j[�@:�i��$���pN�8r'�c��5AV�-�C��v�����uX��@R2Wڬ_�%ӭ)$m��s���Nw���[��QUR^t�c�����H�f8WU%.̋�K�(~i8R�\8��ӍV83G�J{�
O�l�%_�˭2r�����2� T�℻C0/K�0_�AB�#ol2"�AJc~%�Wa��>��e�:þ�!*����q��r.��A�S�MƉ�F2��C-�Lӈ"����� W��:���M+B���aĭ��C�/��Ɖq3�!_&X����/b�[J'ӡn��8�1�4M��9v(��p�)��7<�ؚzP|������.�4���ͫvYy��L���|�Ǆ���P�|���Բ�5N0d�^qx &�S+c�عu𝚅��-$�@�L�msP@�B0�yM����B�@�т:�Rt�����h�����H<ul��u��{�Ot�LV�4N�]��� ��5&��)���N����!�I���� ��<�܇ǹk|�/�Ϛv7g#�?�\��>�~����)r��Du���?����i:|mA�����zD"��P >��J݃T��$���.K�cT>6��[�˾�e��a�f+΁ ��&�z�8�_�'.��|�S�Wˣ��� ��v�yL ��`��,T���j]�E���2�m�`�,M)l�2�"S����$s�#3یmd���	����H�9K��W|�HU~�9��Hdp���j���$�ۃN�J	�;�n��px"CL���?�W-�TY����K��
�b1��!s��P�Q]|�g����4�������ߨ_N���v��@?����B�d۽ʑE���qK��~�Ԙ�@��d�o��z��w�qGYŧ҇K��+]\<^�Ju}�_�Kq��f:��a�]>����h�M�3I��S�j��5yqT5�����n���*+jX�s?�$>���ʧ�����En� ��7 	��'�� (O25�G��D���"��B�(�}&�|�&\�%���:�#d<�������)J	p�r�� &��D�ϩup�Yw�Ͼ�7`�	�<h��U����|kE�����n�JS��\�Ž�5��ڝޣ��33j�=!s/���dױ���Wf��[*��@&�Yv`~/�xccu�i.�Br��Å��Aܪ�2��]R'-B�;ȴ����� ���Ѯ��1��,�md�6�;���m��!�.�en�Ag\��1i${7�G�q����m� ���(o��Z�}[�{;`Ѱ�rle�*�er2���52�_�Xpz4��+c�ud�2F�s��	X�64�l�P�_+"'�5�eY����`rE��s=� ����� ��z�8Y7QG) �+z0T9�uƎ�jq;抔)M��u���_�Z����yْA7و4����S�LCQߴRY�d@��ށ��R��;�׈�H(�J��5G��	��h�_�E����y��DACr"�֧�ֶ .��-ƆPD���s	���dC4�v%�O�����[r�H�!�a��g>3��!FCv���S�j�`]�fy�;w��¶�bi����hiᡴ�=�`w�b���$�?|��6S�<g� �ũ���P�/�ۭ��D��'#���[��b�E���\�$
qo'��'�e��h�=?���b�E��'.ƈI:GS&�ˬrxM�FX'Y`Hl�]���	�
ʴW^%�=�m��Rv4#T��̶�P5��������~ߝ�3�'�������$#�hk�����kNH<+aX�6���&<o�*¯���
�ƴ�����96$����W��o��=�/�ʟ����<��6���e�R����O��EM�z챸�dy]U�27%!�����Jx�/�|���FI�4K��d��)!��f�t�jA}�(U���^�%w�2�>�W��o�fa�
e�;p}��iE.�U3KHo
[řO����Xk�F���.��]�
a8@�����)��}E���w"(�����Wv/�E2D����?q2&ՌIS��?�OU�i��*D���?�-H:�5�v��;b�ko�KE@ S�؃&���.x�[LNoVL�շ�f
XHِa{9��1�+wkuh)�S�*%�5>0S�=;u��[�L��!)P�,����Nr�N� �Ҙٙ!�v�A@v�`���ݕU��kf+7�.����Zsޜ��SϏ��Q��]�4�,�7��A5�Ĳ$���lԼ^�	��:K�|8qz�A�DL������@+C��:B��Ď���|��R���ݛ��3�)"2!H#iu�՛����;s�<�)z��b�QߧK��I�Jrz_�'��9ʏ�<��K�ּLq��I�Z�VMŀߧB���_z�^���n�4�i*��Ea��.�s�Q�h�[���-^�Dnh��A!��S)��MnG\l���i/��=�m�������$k���col[=��F!����5�C)���A���ܪ�:�2���{ �}aŌzr3�F�m4�?2s��� �ͭNƀ7j2ӗғ�`Ah����5�����B��{QY8�A�W�y������j����a�Q?빬��1�k)�{�a#�e�Y����_WS�� ���}C��;Q�=2���Y��ͨE,����ߠ�/��ż�C�O�KM�h>iq�{��ԕ��u�U��W�I2�ﮒ��V�Cب�n��T����7ѫ�n]N������t�XL�J�#����%������.�s���?��Ϩ��k�se+���cGj���U������U����:��	����'�݇�zfHN��|�s����C�4�Q�08�������L�m(4O��Px�s��Og�M����;��� XA3�f0�Z17I�q���j�Gӟ��2t������UiG<�^���*�K�D>ذ`Ě���C*�sX+����p���e
����vJ�N���$�bcA!,4���R�� �8"�~0��\����h�g������\�aa����(����iߕXU�:<ص�N� fT�d��3B�Bbp#��"��A^Pڝ/�M�:q"]�� ���wäo�!Y�`�=�����pI�d�?��Wڣ�}��P��Ё�ρ�E8-~ShZ=ѥ�D��������"�I�G��q��"t.�8�;���e��c2�y ���5��Q|�׍qS�����.�������;�?��y��,}1��f��c��v��(�oS��R�p���k۪2)]� z�)v,U��:��WW�!H�5�``����O��c��ٳО'��7�^Cn��h��(� rVv�5��|���-�?*� �3�
d�u�x���M�)�̈́8�`�N;����do0�Y�)�+s6?�ݘ��	�b��{/JՃ��r���΂��'�0[��x��%q��t�Y�2xMf�l�/s{ٴ�]m@?�[Y���S�!���H�p?�ǘ�!^����|��E�<tA��fɢZ�/]橶�;7M���@Ű2���哖>�f�N=�p��&�����,��l��������4�]<���[&�T:Yd(��i�hG^!`U��h�?~{DJ+�7��2
y|*I3Z3�I��٨ miȩ�Nr�dv�S���}���	��{d�xcX٤!��i^���DT��T��RÎ1���)�xS
�s�����.@X��͐�ٚ�#)��ٷ-�.��93���S3���3��]R�h8h,�B��K{19��Gз�pree���� �̓���ֻu>{"n�\gD�G��06�z%�Ŧ�	·��$*�D��.���b����3���#o�f��/��v�����;���OK/���y�h�C�QW�!|�dzܥ�r`=\f%p�M>Lu��]|uf�9��2�";җ��k��;� 1I��]k�%�@�R2�ZZ�{s%��솎�A'���?K�x����V���r$[���pM	5xn��C��rªL0H��n6�<�P�j��CO_d����M9r-����k�/�����U�pI���w1�n�%�uT�(*1��rج�=�(�In���-�t	�2�;����^%1�������c@m��)�D���X�����D^���F���!s_�'��,�.1�r4.��`H/����\PV�7:���k#�����e�iC��x��uC�Ӎ�
����F��nrT�5�[�Q�j��,w��]A.uQ��;)�)�K%�cB(��� Ow黳X�j�w����I��gh.��i�68�<]����٩J!sx��ia��)�^�Ay?
>m�k�:g�G+! �FH�h�b���0��O
�_��f�RqY�{ɝr�V"�@*�P��Wm�^�&�Q|�1�9� �s��:�U�Z6��@Q��X;s��%:�l�4�e�%(�z;���R��`HD!��g�!k۞q����e���9����}6��eaj����Y�e�l�8�e"�r*�;Ư_�#5�8e�5�H��r,K��E
yǱa�l6�\�\䞰���{ }U�|\�/X�N���V����6A־����:ƀd\�?ݬUb�)�K,ӿ9V�h�n���E!\�:F���JU�ߌ�;&D6ʁ��O��_b�<�_�-A6��a��Ԏ�`%�~L�D��܁+�������ȟ�Q�s*%�R�
�V'�>�6�r�A?�?"�JF1o�#�H��ӟwO�e�m���)�:A�7��������NvɚA��6�g��i��~�w2=�2�݊��v��冸��jf2j���Kc�i�\F��އ�Õ���Ͷ��@�e&I�~���&�����"�z���h̖[����r"��v�-��k6H��������4]�X�u<�2���9|I���,���,��Ff�+�N��i����w88룿1��wBg�h�ê�җUh�x��*��[
�=Z��ӂ����~WV�~uIPW��ohUMo�����B��w|Gɫ&����Vw����80_����c�+�G���M�%��kn�
��C%)	W�~��>�/���h�z��n�~���Y��A�F�7��U5+�wO�R�GhU�Td�28��/�s�%ix�_FX��ﵩ=�*"�7�:���"t_�D���L`�����1��N�X������;�c����R�*߲�x\j&���ęN^�/J'�!_�u'�����O����p�j����u�.&be]&�U��:@,�S��iB���i	++>~������
��Ż�V�z�O=ޮ�;�Z���Y�p8��`-UU�@z���V���&�0h�2�N]�>(�<`�����V�ϥ�i^�Vџ�������?�o�"�P��9h�4=�E8���#ab�P?��Ѐ�������	�l�&
����r��SL�vo�L>�t�����(��wD��yE�`�J����p�8����0^Q����_���t��\	PM��r�����ń��MI
l�e`9R30���R"�3����Wİ)���ˈ�L��p�x�^�w�?<��w���4���W�ś�P��������&�7)dj��!"b1v�� 9�"���4��='|���T�\#�?�R~Fd`dVA�|F�~���"���-�W�� Kf:���kc;��#�Ȃ����
��K]�F1����5�y8�vi��D&����q��F���uZ���N�|'���.v"1����b��@k}x�6%��6��W���Ҳ�0r.5�z;�����KO�v�RA�>H���l@��X�:�Yhq��\�M;S'�3��l� o��tc��π"Th��_����k����^T�P�@���p|��E�T0)o��ݨ˾ؓ��������.�=�6�t2����Yn�Q��e}��X�-Rd�d3)ZL͇g{I��J@4�J^ y���S0�`9��J=y��Ayn�&�$R����u����RM�)j'��V�>E�	��� D��%���F��l�$��m:2�^��I,T��9�=�� � ��d�@S�{O���
7�:���>��^��-0�&�u�������z��Q���r�Z�x ����j�x9۬�};��w=���RL�Vň0p���չB<���<\NzT|S���F7]{ҡ�d�A�q�%}�l�཮�W�0F�*�������M�A�mԣ���F�����r�k�'~��y���+R�J��?��G=0mV�ޱ38�r+m�V_Ŏ˄[�S����L�A�ӆ��������xmf��˕ҾR?dzI7h��y�X]v,Z(%`�(^'5W���J����8�'@]�VcP��HٻR6���Cy�l��dr�甥�F���8�;?e��w|���5l��"�����H���v�>R�)���|��S ���2�_��]�٘{Gk][��E�o�AʜeiŅ�v�)��-� 6�!���4CͶ��V��̲LY��ś��C��"�I���ַSkG<gk��(��hl���u��F���@�\p��~=7�Dprar�U�e����<�pvq2�<�k�kC_5*���-<3��&c����S[u,[F^/?\���=����q��o-E���a�QA���ŀn�KJn��pN�ϕj-0��潄"���
3�"��4pH���)�߾l4�F(�9�&�ԅ@u�#p�i��_d?K���!H�*���+��Y�$��B@��$	��za����Jh�lx��#�4)��xl�{D�f��B�
#��rf�8�ܹ�b�^/�8bv��M�hΙ��\�"�3��M�{F�D�֌�vn�C1Y��6!)�1MZ�w�<Jb� ۙ	��H��ڦG#��d�7�.��rFtmoRGpr��r	��qΑ
a�1h���_���¡�x�w}.s�f�`���I��΢`���Qgp��']�d!v_�79��RU�چ`�T���3��R�4ڏ����s�� ����
������&���3A���נS��
���Ơ��U�q��w��pm�<\��H�^9�� ��wg��Q�'HMB�Hz�8:)�T�`: �;q1*�x�O�[��eWzB��o�v^�	?*��zfݜ������a&�>G~�����UM�h�~�����$&-�����B�.>6]ؘOT������:ͽ�]�R�x���e�I��I�C��r�s��3����{&K��a0-�	_G����Q���rNJ͞x��1��<�Y1�>si����b��"�E3oG� d?�'O�%`�����6A���r���ȗ�x�W�	C-�2Q.��]ƌ�9�2P����S?ɖf�-?xC��u%o&���@+ u��#���wEL=Cr�h�+��w�I�-��h1:?��hi�?ТM����J�!�,:]��j z��%:����`!�17��������{ا��(U�c��G̕��e%m�Y�[H�`�G��8S���Τ�2h��'γ]�|7�ؐ�'SCO!r�� |f6-J�}���;P�4����f�_�Eeص���H�[P��Gߡ�<�f��Ǉ(���/��P��#����_�m�"��;V=����f�Ǐ��\v�I����-�c�8�������V����>�>��`l%�V7w�m�^�Y�I��-o�ZP�v�;���/��I`Ҟ�ߚ�<��؇_>�'`�[�8���S�S�jW4U��4/�����b�{X?�ɥ���T��l��e��ăeE)�"�N`�Ϟ������f�?��ʏ����^[�/�E�W>iZ�Ə�sn��U/��RN��ꈿ�s�񟘹�tYxh�6|h�^@�Ŏ}P.S��Œ��Щ��J�}��QB^�2��� p���=r��8��o�u���yx�_M�p��%~'甃�+��vBI�J��Z=5�,���ڳ�Q"M��=�AU@�����r1�tܕ��G^��h��R`,�X����pС�f)[�2{�x�A��^?>��bpv�a���cH��:�%�`�X�f���tN�r��vFJ��NVj#���s��JL��?�1�ͬ
�3��N��9J�\���YJ���у��@���G\x��v��ϗ�q��)[<:1���4q-ߢ��l/��nZJ�I�*ľ�@=��Bs��J�ʲ����+?n�C�e� ��l2��@bp׭�{9B-!��1���t7�	g�5�c.T��^�0���E���5���x\��)w�`��q�R�Nm���'_�4R��3oc~�XZz�kH��y�m�"*�gD�I�'n�GԮ��b�	��c�)6ÞM%;~R�3\��fz.���Co��@U��E����$�=�(^ߪ2 �ڀ�����JiVV*S8*RSt�mM��"�=Z{"o���=
ͮ�NL��1)�}}f~�;�v�m�ʁ����?���s�FE+1u���l%6���+� h�S���L�w�' ,��'���EM��"�ً�?製�������ĬFh#�I��#\�)U�P$���ea̶�T���M/�dC�Ej�?a�ˎ�ZYQ�!�2��Δl|�58J����3OVU��=�X|���U�o�DZ�+;���ֻ�Yg�`�,��W5�� �@��*)�M�׸�d)ވ�ƋG�!bW��2�[�y���7��2S)�daإ=|��< ��qh����@o(�o� �?�J9��h)*��6�U��z͛����m\�&����ǘ�	�y0��ﭣe$�/��1�������8oC\߯`ܪ�U]2�5��n��M��A]�A�t�I� z<3(�#�����T7����e�Zf�L�bq�^F���bX]��yLj����X�d�3$7-�
�T�"%���a����n͹�;�n�(A���V�r8�vJ���Ez���Cp�G*B5�o���a�m����f�������^RTU���vo�r0OyO�-�Lx}�쐦t�]+��d�	4�%27o�V���y�?����e��V�ŷ���~�i�1�=`�Y֑�^�1m�@�z
C~��ϱg.\a�G�$��#��qX��=�����u��r�jf=�!���gZ�3����*�S�p46s�F��-D|�I��D��!n�*Ff����CT#.�~�Ӳ�'w$�N��������#{�}F�!��o�|��ҷ-��� ��m�.�6T��PG�M�P���7����A�4?�pV˿��%��k�<���]�N�s ��!+��zv�DO+f.��B?�waR{��h�XD"ǆ����7�"A��%�ʐu�X��t�VL��J�:�q�\�A�0@DD3}�De��U0tp�*zv�W�p��ibb�*J�>K�� �a��{���Y��O+m�3�v����3�Ӝ 8D�N����ms=�e~��J�MS�F�{��HC�3� �rDs��T�!`>�N�"p�1;j�?[a5���|nwD���$�-��h/ʳ�R4b^lV"k�;��!��k��
�1~�>!֌6�rM�v�jg���E�0=G���^�N�>�l�.�1�DkVd�*�"�H��DP:=���G��TA<��?l|mR.���(�Isޠ���l���Z%��C/E�,����QS�K�#ha��G\Q�� �k�O�%��N�h�Sy�3����{�
����w�PK���4��&E�"Ȳ=�AoAH֐�J1��[�s=���n�K�V��F"�O��oW��&��i|0{�4�G�����B<�5�|�okmJ�� �So�eK*�5��M\������M�ےS[�h����@A��5��!���"ٲ�Nwy��|H��:�Y�$	Uyni�<>��Z�b����<�@�l{9�|�jo�1�p_�=:'��EC\=#@!���t�����)d��RȬ>>��k@�W.P�MԌ�t���7FOأ�\��X�(���x\�ԓ�ת�l2�*
��.W����.��k��t:iGjC����L�ǉ����;�׫���
��ҫz�$�%9d�����WJ�K����GY`Q��X���D	��E�f#jU�& ��`b������bh/_r/آ'���|�5HF�2�Em���*�f��x���oB`Q|,D�z
1/�1��!e�P#Ԋ�Ô�?"z��(�@;��M�h��]�d�4W&������n(����.tI�/R���z�Ѵ�˭��Ȕ�e���	[�,W,z�`����s=F�0����߳*W�1�۾J�r��5�pD�n�Y�ˈ�n�u◧��Êm�I���?�YB� .��[��z�+�!"���h=�5j���R�A}쮽��,P9;Z:k�3��P�g���T[���҆�~B�q9Qij��nF2N�|�������?'K�O��	F�����9�#ȯǱ|��T�)��7�u�xb���X?j��*gB�r;W���׫�4H*�p��ų0��Oo���:�$W���^�a������O�(씂�;
�Q��:M㿙
q��P�p��7�B����w�9&��T^��}4��b��"�ِ#�G���	�M�uS.��j�@����E|�J�]�yEw�vz�"�w�{�� '�� �u����@��,��Kȴ�;���^0�-��="�����pjW���#J�*�#����yF�����DNՂ�'i�X=��Z��uj��5Z�2�ʰhEN�~��R,��x~ȕ3~��F��Ê咓oopm�L��οը�Ze���D�����2������b����߰��@�=+m�'�a�8��M���;w"`F�A2,�.�L�B�THu �)Z�k�� 9�L*�Ԩ�!y?z4Ή��f>`\H��B�MM-�yY�h辵�Y�,���UL���t�A�dӍS���C�:��8[OeX3�PҔ�C��ο�:һ�6�^�F:$�sQO�b��J�7�'�DKx�.����%_����BŸ�(K'���u9����s8>U���$��[l:΂��F+a����i}������N��_'�?0<s�m�㋐#�%��n���s�tt�sۆ���Ʊ��f���h��P�2��xFF=���8��=XUPCM�7��E,\�Fe8�ƏI�l�Q�K���i��1�P��Y�G7g��UEn�ٿu�}��;������� ������L�@�����H�j�l�4��s���Ȅ�^��[@u`���ܭ�j:���t���������U���5H� �S�����&-k;|�:��=YHR(��bӐ�G�. �rU+5-�T$���f�����T(�����?h��-;&pC�+���+߲.��lg�_������ʳR�� �U�GXѯz�������y�ڧ�v�r�8kk׆(��glM�MH��<G?i@�98��k�ሽ?�x�K���=���5������ߏ�(�)�"��; �]����,]WC��=!�(w	+8�B��7_K����y��z@�U���-��>�t��y �H�37�fZ����Q�:h��G;����/N��U�\*[�����X�J��
�у{i}��7߶����̌��l������c@��&9'�����ӏ!�'HT�Q���85:�G���Ā�kݤ�ő$U��U�N���]-|m �/Ӛ"���R�';1FVسs`.�b$�'3�~��V�� ��âe[��(�V��4ŵ�v�|>(ŝ+.��5 ��m�|�l�ֹBJ<(��fy�(��%C��f��$WIe�i��0G��I�����TG�2a��9ڍ�%�!ĩ%gA��g�h�QR2�2�6��隱}.�;r*�9zҢe����>%WJd�yt5��T ���RL����6!{�X�#+��K��8FƳ��?\�9�|\�t����?%���� w�J�0P��f�8y�l <>�ߴ��ܻ��p$g���ϐn���C���*��E� 6��nXbw� �f�LWR�ee5�rw��Fʓ��yu�������؈uFR7���%^s���B���t��eu��M�nT4�K!Vv�b���r��d�#@1��> I��HpA�܃)�7���-v�I�8S  ۘS�E-c:����@��dM�P��Nb�ժ]���D�Ű��V��`���eAa�H�:���Uf�)�*	�"؃q�2�~~���I6W
U��F�f�囃ls߸�3���Ԛ�p�KPG���I��/�(g�  ֩�����c�l�D����Rg���&�����X�K+:��o��T���c�D�����6�+{�YW���Y4��D����nCGΧ�u�X�lS���|'�'�	���ǘ�����J�JW&��ZI�c��y_��9��B*��qN:X�odj9�%�c�ff��`T��d�[Mh��x����l(����Ff0�]9�-@�yG~����.<v	�$p��Qf$��XC��t�A�.rYt����P��"XP����S��9T�C��$��>�nFX�A�i�;d�$��U�����B��|��|؁r�k۹�&�N7ծ������^�jtô�� ����M��jKk�=��xp��X z� �������8U:"�F��.o��#h�3wm�t&���%���������ȓ}�YQ�	����,����s�0R�ܓ�/��\��4��=��н�ډ��6�
W{3���f8r���ޤ��a�3�T�d/m/��]F\<�,K�m��DShS����p8�{�tѻ6O6�!�Ѷi4����Lpz��H$h�iu.����*����	�;��8�_���N������mZ;�4j(%��ȅ�&��{&Z���|��r�ne3l
���If�U;b���H�ݽv��+R�7�KҾ!M�8>K4��dW�G�*��B���3Q�g�F��b� ދC�}���K�b���H\�[�a�O�v�ڲg!�������Foډ	d�Y�� ��l7y__9zH���� �7q��	�b�[�2I�V"��[	A�d��>�jT�h�]q�M�5+(=O�q*���o"���Jk��IK\����C �)����~�ՁT@��a�����Y{L�O@n!R�ߵC����HY|��,�ǯe�:���������{���Y:]4�&䠧�ԙ� �< N��7��CR��w7ox�p��"\F�D�!R�f.��*}�?��u�i��4�e���k�uHI���ӷ�'gJ�g�3J�Vd��e�煠�@	%�}.;������p�����蹋�n��Q��P�95��M~���D�[ұ�uԟ�D2�+eU�r�O����(�A��(���V������I�
�*��qV��r�϶���z�� e��3�1�.�~���1x��b�@������E��:J
y��h"��Q�X����<� ^�@~2�����.��xٌD���rE`%��H���'i��4�=�J���_��42:��{9�x�;�BK�[L�!z�� �Q��!lh�r�o����M+j#���s�\]��y��"rv�
(��E�ߪlcc�pZvQL�!ddX�et��~.�زP�m5႙�O���7:ݏ~Ž�f9��@Zҍ%�w�F�4��c�M��}R[ʉ���G��B�������E����Q�7h�T��tj����FZ��BX����P�"�e�c����=���^T!��i#q/���D����;/�\�D���ْ&j�(D�|9Z�c�����=
�����rp�J��s�a�K�x��d���}�~���F��?�|�v0��LI��r�	��3���|2,x)��]f�G3-*d�&��ǜ�!13WPp^�F����in�t����d�tbC����o�հ~ْZ-�f�m�t��	Yml6�VX�,�׃����v���=(��ǚbS�P��p��Da״S�
�쪫�x�RjB.� .�H�JW䪎�3fx��{���`^n5�r�Ώa��_��[��T�޸d�*+�7d����.�AqT��(�pc��Pp���^~���<[��%2����J�[$V���ñfp����5�[
$��70�[�U�z��i��]�D�4>�e����� ���M�T_�� ��D�̄A���#J�B�~���*�1p_�A��B�o��E"����'}�"�/?$���
2�mjmf�]5����~d�v6u�z�T-��(K����g_�ַs�L�+�b� |�$�$��5��0��5�n0Sl�G�g�=�#$_���$7�̑+�CG���vå����q�����˓CӨ�����S�,&���V���_�
�)k*6�Q����3g �����XE�}n�pj�D�C|�N� ���J����n��V�9��l��>�
����T��NX
a�@D�X��\���-0��E��0p#����*Xl�,ifm��Xz�-� -H��:�ܗ�u ���Bי�p�C8 ���* F�.����25c싊Y�q'���l��_9��X�vĸ��� ��F�gK�D�A�!��(]Y��V-<�)��2�Dn�d":S�]�8a�P �,�L��k�����k��8�쬕��S��/�*��L�@h� {�Q>���Z�?"Rx��C"�7��hsPc9����Z�`X��Dۑ^�����NB�i��, !SԯgdL�B�=!d�0-/�N+�7�rA��(;������ҕ�![m��V��傛���A��OMi�(��;>b�V���c.L��D��H���v ����(���Y�����%�6]d�=�NL�9�.�S�3X@�I�a��ZӷW똤
*;�4��[�7��_�>�MP�,�����߾���v�#S�6;�w��
����LF̃�3�O&�%5��p��:�ӡC��Hˊ"�od�'29H�U�����af��Љ������R$��E����QC\��s6�D�t�|Ό� �4S�B��&���1�ʌ8Ҫ�l+�x3;=���(�Sƒ(d`����%���^j���/�je'��-�2����_
�;&9�EA��~��e�W�Ը�E𠷟����z�
.Њ���Q���zܗj}�X�7��ۺ�X��ܩ5'��k���r�����ʡ�#�.z��-�/��>
j}8�u�<먯�t���U&m�Ҏi�>�\�I9rH��"��<�|J��f$!$�Sgt���=]Η	�F�K�.�����\n�+�y_}>����A�M&�����w",`�Fyx��F
޴y;S���Qd�/Q[�qo�N=̽C���m��M�W�Dqqzq='�x�C.g��\���.�茽������s�|[ѷ��L�����L1�{��E�}�C]0�������Fwh��r��8L/�R��Y�����!�_R��Xҵ��F�#��E��MK�>+�r���a�2��fZ;E&��P��Í�P	�D e����u<�cGЊ�f҉ �P9��gb'������(?c`V��.�)s4�%�2tl�Ej��ew����b(����X�ޒ	��Dw�I�_Vߜ�����0������TF��jK�r�f�>ͭ���d�D�l�S*��gO9)��s�,�J�u�Ī������r#�Ґ8��f���e$<��%+���e(�Q��è�hE r�[�Xi��Y7̰gR�m�h�q�~a�N���.�Njm�ǃF�}ju
�� .q�cVՒ��4Y�LG�65�V���}�r�n���E}a�2>����D�-l��sN�d���Ց��6Ϫ�]6��R\׼�`�Ε�ATˎ`�D���Ǳ&�4Y��l� fF����臅ɶ�<o��V�
��:�����J�<��QT������$�O+�m��m��\6�F�x���7z�����"��ԕ�?1�E�v}�%榏]�v�ۉ����ip썔�l���h�(�>�k��V�zL��L��<Ғw��Q��]�P:Վ�E���@�scC)��wb�GvԼ��5>���d�tXn�S��q[���^{����	�w��e�u�g�v��jgp��������H��M��}Uuոծ.I�V7x�N�E8�I�w[o�G*��*�s��Aм�7�6qߛ���b3���ٷ�V�e�P�<]�͟]g��`?�>�P�dQ=��q�y�3�a?�tF!V�G�c�ʊ�2��{̱Ҍ
L���ª��z��X���,A/�������p
���(���!�7>�p_Vx�l�/����.?��
��@o]x�[�
��>,��� 2�2�a���O��c���oi���3pVƗ��)�|�N?�h|���,�'�����l��vh��Z���eiM�������S���+��q�|���D�~5A��~vn�ӹ�ޙ��@�7�d��!��z`�t�S&�b��Ku��	F%s�ޗKC����Pk�
��j��;wE�R'E�k� |�����f�Q�Cߺ[b\��hRn�o�gVC^*$��Fv�/��ٙVJs��k�䄋��j�!��^��#�2��"��W�9?�W*�3s=+zk�� ��7V�i�nC��8�H������s��/�]����m�S=�O	n+�Nu<2�WM��^��	�$�Mj)6�0�L���8�۟[�a�<b���To#�e3y��A|U>�T���8�53T���5�u(o�r>�و�IѪ������c��l�$�+i�E/[T�%&��7�����q��x-�r
�;j	��.56�qTtf5���W�$n��k]d	�p6���u�D7�3 ��t���`�'�2A�i9��yE�OJo+ԖnT�T�:�v�^��}�{8rV�2US��W���0T�z�(�r��1�HM>�_�0�lr�14=�u�� �?mZ��~M+�	o����Y��l���=p��,Ԍ��"��7�T(�P>��_�6w�m����ixg��٧q� L�x�ZC�n������ O���y�:�yq�B�����&ŗ�OS���O���Z�f�dM�w��ɡ~9Z���?���������"`v<%v��3Gn���+�g��H4;=�1�Ĳ�'8�i{�O��e��qH�S}^R�!�X���R̽-�oY��?6v-L��w�]�y`i|����	�LZ�1#��)�����G��JS[��X:���5 �ׂ�ŅB,� I��D�~5]`C�L2����~Z;8-��2=�����WQkRU����/�����v�]���]���_���`m�*��4=��g������_�q�vU�GHj��lA �r������XKM��]m����s4�Ȓ�<P�T�5�We"�՗k�0���i��ܺo�>����Q�����������{��.�)�$.�f��O��X��E�;P	1	�v�y���)xs�g]M ��r���J�m��ocF�B���gAL�PS�hi;C�1��ޱ����@��!�1�����C p!�����O�#\�ȨVv�e��Zf����-%\��)�P�R\�W�6C�B�ꛧs�O�>,�{7�1o`�?醺Q�
��N$��@/	]�Á�	|���Q!7�fw�p��b�?%9.��,2��I/T�(+?����l�A���:}3����iVl�>�եf�%��3D���s�B?���b�p�l�������Q=�n!�UP�^MN,eŘ��q�� ?A�	�H�a>7��Ā���ӯ��Kw�_w��Fy)�Hki�`��K�H E��(�����_�}�X�k��^-8���頹��K��D�;)�\>�?��&t3���CRQ��9VI[��5;X Գ�!��,�_�``���D2^�YO]��,|Kè��]�]�L��u�j*�������g/KX �w�Bn���'��[��F���/��VB��T��r��n�:5K�`6��x���"fvB�E��n�J��X,��O?"Pb�|���, 1��t���0w�]3WIl07��Qs��!���ؖ��8�eg��o�@=l�4Y8��_ѝ!�b�t%ߧY��4�L{��h�%���joh���-��kZ(��H���UP�N3�z���xUk��
Q}���g�O%�y�����G���*�l{Z�C�20�y|B��Dv;�[��1�GcM��#9�F��$�8:SU����V��h�\L�X�n�B�o$���!G��>����*" ��M�8g	2�Ԅ�T�!��m��@
9>�Ի�R���|��?O��.Fc��~o1kd���-��;��j�&��+���iK���K?�xS��TB��B�֚�����9<e3w�h�����~�"m��!T󠞢#LJۮ�UwX)$��i*�U�;��;?rB�#�x��%4�-��t"�Q3fa�M��+�-��]�L;����]�{���A�ŵ�}��ʭ�G��[i�������:m��9�]0�d;	 q�ܮ��E���j|^�i���M���b������˂�~���.ˋ�� ��s#�����Z�_�4]�����(#H�S�_F��/�$����!���&Ol�K�A,I(�s�Pe0���#IP�	��O���j
hU�W�wq�Q��
�A��۔��.�aP�`�OP����(����#�9D,ߞ^h�1@�;}t[,�P��������@55�iꏾ|����x�Nx^b�_2��f�o"�z�U��/�����I��3�р1�	_ �	���}��#G��D����4�kB�D�ZH���h��)2�D㺵�;ps���,�'���H����Oc�VF��m��C�	��� ��N�xD�)i��H���ݞ+��ߕF�����T� ��\v��A;��[���H%��|C�S�� \�:�c�?o�	�K �{!��Piº�m"]A�w�	Bܗ����<|Q�	ߨ?C�y�V믃�?��ђ`�3���~R[Sq���W����b9UU�2���&�l��嗴�F�q����������I_�|�٥S�l��Am$T��6Y��q$���X}������k�D��R_���@�=����p%��-b")%V�Z�_�������'���S�/�S��g��3�Ю����������Jv���"{%��8":uƳ�{!�RRj](d��i�zs��F��f�[�����!�	`�,��k�z�X���]�+�b-Ys\d�Z�������
�˺,(yř�͊9S��q��w�X�Y*WҔ��e�-�T�)���H���$n����F�+2�|߉�w!�H6��/����m!C��Vz��:�$�;�c��
��NuPj��k*�l��PdMrC�Lr8��|�EH��,䩄Ɍ��1f�6�j�i��s©�%�1`N�M��K�j���3�+O췩�d큨�.���j�y1�8a| `��5��t��;��ͱ�R�#��o�D�я%�2�xې��T$�פ��i�Ehq]q�P�̩ۘ+���#4���~h�s3�ju�C3;u:͵�M�<R!)��Ep%�C�E�gZ�=U1$�� B4M�)��S����Y���",-o=�?�"�=k��f��<����2��j�F���p���rWOAJ6��Nm��a�SXݱ���]�܈D����lf/�Nb�Jp���s�O|�*U�.\��Oݼa�+��P���E��l;5f�Ӂ����y�W	Ь�v@N�=4�+<��ɞ�n�#u	�9��`��W'�~�]p�+�<1J�����ր���s�Y��@�+V{���mX(=�zzz>)H3���F{��n[�Q����-�tG3�8��RʧR�4��æ��7ħ�g�8��*U��w��� *��cY,7���j�(������,H-d� �t,q�H�-�WH|}��cơFM�?�B
��Ù���f|=R�Mf�蛶ïzö�(ӥ��!:���)R�a�����y;=컓�3�x@Y�&���29��^\���f�~�D�!?}�*F�595�*����F��L;>P��e1>h���n"���<﹦�<|��PY�е��AJ�!�?iۮt#�V���p��߅���<;���3!"��"�%f�a�=۩_�mz{8���[�fB�)�E h\S�zj�6�`�!X�Y/�~�I.a�����ͧ�������:�G4�2V�NX���u���N`/D넪9sV��D��~��6y.�t8�~�p�	S&�`+A�����B�rh|*��=�2���s^�s;�&q¡��miuՄ��l�-k��� �7le��7��ؤ�1BU%*m��>�G���-1��H5���ׂW�T�$^�+�XLڞ������r�竢c�xq���5��ǡSgS���� ����0[dV��TR��j�x���!M�0�g;s�4�KE�����k�����uϼ^�q-�T����?^'�=��oD)w���n�R��P/H���Z�;M=�T���-��P:�ߕf�({g��4Aj��R�v�B��z��lN��q���`A�(6��Ǣ�R`\�����^b$yco�z���b��ԃ`*EI�ĳ��_�8��"�S�t�l�_���^��CܾK�R����S��J�R쉯��:q1G����~���my��s�ˋ�-�Y���ឺ�
Vq�]��6i4�r�!�ir&7o��<����-_؝�����v7�''r�՜8#r�l߿�)��0�ӊc�]0_��v��P��h�B��j��Q�'2���d �˝�Νąq�q����P=�J*) �E�ֹY��e���@K�Λ{ӑ��׈o�p�wX�������G|��s�2�C�W��aO��Ȧ�B��8���O��a�9��z�PN	6�X;L��&�\Y|O�d��8rռD(����<ys�#4���Mw+�=]�(B�*an��8&5��PM"B�&7�A8���u�k�<"��Ȏ�^�.a���0��1����0�V�E�21�^����Fء�W=��v9���������K��[D���4��Y:3��0h�[d��5�(�	��Jwp_o�.gE�X�֪��V�Oȿl]�!(�+I>��7Sc��A�Z�3Q=�o�8�*�ZK���j�/�������h�� �s*Ӈ���lI�����L����
$�_��O?����ꀲ�j��|���rā�z�m�d:��+�F�\�_2�4;�>į��Հ�D���slc�sl�A.����j�{�a�W�-�;,��4Z�F"cU�F�"�*�;��\��l���R�i����U`���2!Z�����Z�b;n���q��r�k�V�s�3�t�.X�l����nV�z��[���2��C7a�w�_Kn=�*��Q�Pώ�q镣'9Z����ˤ�_[��?I�H�,Wm�w�+,�oY�}1��B�IL/�v�Di����z|�yJ��i�t��	�;\��2*F�\�%�M��ĩ�c�<Wy�Q#�'��HY�bEe�ɐ��@��!��'��_(.Xm#! ��*���ji[�#��q�oS��.[�d8� ����CI��_�T	��	7�j��f�KNwN豈��7�!��b�<�� ���=�u�qxU��W�ss�_�@\+b��%�����l��01�7�I�N�o�*���֝[N���H8���)N�>��[9��owS�O������ � ̩eG��*����H��[���'<a�٬t��[%F�3BU6��� ��o�R�-�N�
j�G��OY���/m���b�2�U�~ӡּ�|_|Z5���CR�.0q��q���D,dY�Z,���S�}�M�YO�H>Kl�\(�jA�D��[�4�"��[=�{�5��_��_�ۚZ�M��<�DV����G���� ����]\Ó��5"��T����T���6�Y ��2!�*�s|�b���; U�#����:��RC�ߦ�p�&�8� \�;fi�䲌�ņ�t�rw�/�o�$��t�,�î�8w�[z�Ȧ�[��<��<�I�_���=���K��r��y��"1/�6��ڿ�3�	��R,��c��c�:I��Hsa��AN�د������S�kHb�]�$����܈��ګ�t���AC,�2���l�0��Qh	 �:Rsa+�V6S�W�f�~J5p_���}����m������bxn-�Y��q��3�Ob "�_~-�&k7��#��ƃq�5R"e�؅�-���d�4�y\��~����S�!�j�R���j���U+@kܔ��zvl�M41n��-�헔#�� ��M�草�)�θ�W�����~(x: [J���E��z�?&�uU���� ��3%��%��ֵ��N��r���|�_��\��'3�-	��j��I���g�vTƷ>X���M,b踲��u���j��Tc� >o��N}��>�VP"�4F� ��P�Ĩ߿ߒ���䣪Y����٠~��Dil.�8�a�G{8�p�I�#�i��V�(��:*ʈ+�w%^Wm
`���w�Ջ$�U��}�����{�\���ˬ�t��i�Nh����P$�Z���m!�:��5d͢��'X0)m�&#��0�E������Rb��U>�h2~���#�6w�n��:��l�����W�+��0�Q�` ��o���(�}m�!&M*}��S9�j#�q�qL�%T~�LSbR��1G:���K-�[�1�$��藁=��LIJH���*�7�Ԓ�
�F"'��#��37��4��E���i7�2Pg�_{���-��D�hl4�T��߈�?�@��i0o?.�Y !��5��16�UH��yS���ƶ�6��T��/��	�ǸT���뮶%�g�8G���皢���37G����Y� 3!
рFet�_�jn�;���@.5��)KW+v�>���a+$EC�=S�l,�^�;@�k�9��^��N�����F�\F�9�Y~���7*@Ђ�lBX�0�x�&��{��硢-jH�Z�l>��W�[R!:��ءb��\7s��bV5<C�T��!�a�P|�ȹ�e�ؙ��A�6bc'��=މ�,�����#��A�iu�ĵ��x������e�.B�߅���d@�F�RB/e��x�p��ʀ�u.��|�:L���%�&P�5�?�<-���9�s��JR����I�r}y�f��M�q5��b��NFe������M�\�aԖY/�FT(ֶv���>��ߡq�䞍�����u".�0!��P��P�w��w6��eb6;�I#����k`����#�1��Y֚Vr?�}�ۮ:�pQ҃�ƥC���fKH�#�}�5�C���.z(h& ��c�@�
E��Vp7Бq���0)���%��h�ܝ(/bi϶�'w��CPS\�)�m����PPRZ��D�!��0�I�Kȗ��#�
ZfE'�KMVn'�޹f����݊����ǥ��Y�ܽc*��CL�V ��D�ߩ�7J^e5�G:m���MwC�ko��vA�,��1_V=���-����p��Cd�_��.%�m��g�����򟇩���\�<�6�"ɕ�tI�nN�#��U�f�H��d.�6Q��2\�S햌*�+ϸ>�*N�'�S۸��=�n^���J�r��4�2���#t�&԰�$n�+Y�Q#1��f������_Ɇ:,�H�OǸRW��m��K7���rS?rš%B)@t�E+�ځ+�w�YreJ7��wP��h�_�^6 �&9��%%�
��3xL ��R;B8�E�.��G�@5��b�ϝ����{�no��Y��\!��$_1넟Q��-��ܛk`ݞ�o��x�H,4T�AD[�/�t�qQ34{�=WT��ENQ�[5a��
��=�� g��-�ˡ�)��6��[��Γ�	�mq5�L(��z��cİ�ϝU`$��������I��2H;K���r� ��,�1��v��u���H4+��u�`����Ed�{�=*�Ҡ�����/1�*�	g�<݌3��]����ow5�,�O���q�B����.~,L�e�g�k�`��5#4�00ܺ�k�͞��U��9��b!�6�p	�1Y�ąLCU_��<�6
FৄN�Z�JBv���������g�wS����߻����}�h�刢EgQ�Z���������~$�y�.�8�ώ�`-dj�s�ŗ����ȫ�C7g�FI,�����f	[U:z��{�������˵0'm�wI�
Ȗs�.�F�.dYu�(�-xa�g^d��@����/�\ �+�y4!!��
�d���y�� �.37@~=EF���#�	l�/����+�5��6�Ь�s�1h'Q/-5s�V��H�e�:�%ށ�@[�@l�-R4�3B�r$�����݌O�s�k���I���vڱ~�X���嗓���^Ϋ�f+�?���m����Oݮ�&3�&��B�C�!K�܊EM{��|��%ݷ�)�c�K�)���Rr�w�jyy����	���1#�K�!$?<8x�d���	����z���o�(�\;�bM]A(���J0��S2:t�}%WL���{ݟ�f�fG��z���[�u_�����Z#���']àA0�
�H3�3z�F�j�$շe���\G�W�=����]Iͮ���+cW�`�4"`'�W1��s�0�s$�PE9[�������g¯�����/��4(�	.�]�P�كYpPT�[�@��P�7���ZY�l��+G~ f�i��˛y�T�;������gKT�!6g��=��]9����W��5A<��'B��N��O$�Dq�m�5�3��φ�5��Ƚ�y`#,�����82<�Ty�q��m�b7Ɇ��ɓ�d����?G��6#���%,&�g�Z��|�y /�x��\m'N�I=ay���ll��_���~_����o"����M삆��+�,����F�]p� Ծ����+Џ�z��;�f�SԴ)/��� ���4|NeA���Q�
"]��+ԭ�f]Qʕ&���M9,��zށ�q�E�X��Ɇ�k��8�l������ڟ�Lޑ�����LU#�٠�C��h��E����dmn��I��	�w���/]
s������PcM`��"r^��W�X�4dv��V	��ؙ���čγ�C�pk�����L<�;_��b�q���&����H�b*���R�E���f7{�+/Jeo��/M�О&�I_!"����.r�
7Aͣ�]�z2c�(�~b�c�|�� �B��rk4��`,H��l���դ��Û!+`��xJ�V�§�WƲհ�=,B2XYe��F="�٩��=���˙�^��I��C�ʅ&������?��b	��Q��zY�q\�g�m��e�J��2��P�!�FZy�p���@���g�.Cy�,sE��O���f7G��W{a�N�L9aqZL�U�� �A�V���ût�J��W�����~��f^�9���P�� FO&��;Y�bv��o5�c�w�v�(U\9�k�}ݒ� �cvQv�m���b5�oҿ�S�+�oC��d	nG��D�)Jl�K�}g�������7׌Q���͈��I��e$�٨>��F���͉?<�7� [��Fi���ř�}��P%a�,۵�m����Ls]#T���_��ݳ�LM����k;Z90������@�=g�^Gؓd1�W�tq��n�7C�q���l�s�d����+>���qޙ^�&��WӶ��"4\��sFj|y(���Vq�s�uıƄ�|X݅�#����PF��2T��b�.5�hR��ʕ��9ȥ7VD6��B�[��6�:}f|!c�32��%$IJ��\5�dm�t����J�?K�8N���	-_j�:���t���Um�X)!�r��3�c��ލ@�0>�3G�_�������F�4��Q�;,,�1�@%&t�����o���l�тd��U1�0��v1,.���/v�_�ag�9d��>����z�X�1������L8���2���fXa�8}@���h��u�G�M'��ج?�Ϗ�i�Ԏ�+�#��z���뙒u+"�h!���h�) �ʓS�ٚ�ڕ�/�����}E+�kG��{��� +y��0A�6[V��m��{����)�$�4�=ׁ���5�bf���z.b<�|.����g${Ic�e�4�����-��u,'��;T 4a՟1��@�?Hr0����b�!�Oafλ,�RS*dA���s�3ޤ�F�ʨ�KP|�t*͐($����Ohx$e�7�~/@��FL�-�A�{�(�!<����$�����=�i�Ol�;��۩e���~��V��*�ϒ'�zz�֒!�.Hw2s��/���_q��U�M8��=�U,v��x=Ѐ�~}hH���ӵé��O�I`3��8u-��䠛���^��	���F�{�r�*%��4s���Õ&rRrf9&�\�12M!14(>W�H�� )��G[r^<+�͒Mf ,#d楉*�d�i��Y���i9�s�Oia��,��U|�f�ՙ�9t29�Ѽ���ErPq�� ��t0x�]�b]F�o`����wVCK1�� �?p��wk}��Wƥ�˘%=�jB>��:F�}�S�#�����'�Ĩ�:�@rp1�^��4@��BE�Z~�o7�F��qxE_W�(-`�S�n`�s2��^>A�1dn�	g��Ӱ] j�����?G�aܺ�> x��WX0A�����ь��f�U5Lo�"�yP;�
F�q�������Ũ�M�d�~�XNZ]����K���<J$���~�F�y����y���#�sP�7���	�s��<@WR����R���3z x�`g$�6���4=������NH��r��5�`�}2����|Yw-�eBQ!�2B�����K���uq���v��ׂ��m2����;��"�}�d��%_��hz����A��7��sS�����n	�#ZR�������#�� ��$���e��j�ij�a$��-(ٯEki�m���j�N�Q�^*�x,i�Y]3B~SP��ʳC�K�K*��,�f�x	{��6/-�
�3e���`�((�^o|B-�u��#��f�y{]�˼2��R���w���Q7�
j�م�Flz��-��W"@�j̢jʙ̥6A��j�;Ҍ>�Y\<P55���g�&l�i�^7yk�A�q����3eF�V�T����!���o�2��ag	BG�a���V��ٞG���T�]�;�n��M��b�o��p��r��6�s��m��gT=-���+wB��	���auN)�Eg/�?�i���U���%�ψ)ك���7��c5��%F^���7D~���I�w�4�W����Ѳfh�[w�n��[�7 ���	�d1H"5`s_��_������>�S���n\�^���\mo	�[�':N=֊9��˅E{w_���������F�5ӻ�Q�?����̒`\0�XR�(2�D~�����uu|�ʂj2~��W��5����Z�z=�F�ƭ�E��l��ð����^R|_��W��9�vL0�_�硲�T��"�6"��<�u%=�8" R"hK-���2{p&sɈ������i��;��m�����&C�@n�)/��\(g$V:N�KɊ&];�Ϭ�	��@YF�5�>!X�Gb����t�������W,W�e�
Ns��6Ox������0L13?�y��*����Aa��Xb�v]�4�kZڳIk��v��V�\֕%ʢ��;z�gL4y^��0���/�ߦ�,�̨��̮��2���*e��0lHoF���������#�����Β`��X"�X̰����R�2C�قPjm׻5�F�\����^Q_�zX�i�υ�V]�h���u����N�-TS^�V�t/&M`l���Ӈ�:6pV�u�'��O� `��)�&G\A�r')���y9U|������%�Y{ņ���.1<��.9}���nY/��o� m�ECN{�������i^�ի)���Ht�y��t��K��lD"`���s5󽥶�LG6U�|6��ۋ�ҷHL\GY�>ř͊��Z�c���������UC� �S�F,(�7�N��	��a�9�8���`)l?"��ʛ�}��_���h]ŧy�Y_��O�$��4�Z?�Ύ��-?�N��^m�m20�1��F���է�!	�u l��T0{�=b�M� +UKE��� ��r�3���#�2�¬o/KY�4�*i)̴�:Q�m�l�0�P�����"�hf
����2Ӫ�iʪ
uOO���<���@����D_�#���,�*o�*w��G��oM�X���\��is�����A�{i�B�(3�ӨS�]Gm�A�u���Y8Q�pr��N�NT�x�8�D��
�c��"G�y2��r�<ke�L�O'ii64�ђ���X� bWB��Sz:�-%f�2�t�D���ߩ}��.�cq��{/�����t|�����[L~�I��`�`��JI������8D��A*4�f{Q�te۝ҕuѲ��
��_�f�ד�6=y��f���Q��H����@��+���uP�=��xz:�����ܤk�����a�o-5DI�*��&�O*�|u5�`F���y�o.z�2��"�����W�b��8e�	�v�U���k ]�[}a�;� �1{����Mdh��G�;X�OF*�l��&%�掍�x�w���2�6�U$6��@�k#	�}RӔ����6S�3��?���P̑��H(�X$d��D.��� ����k�V�^?�&����][���y=f�+N#������W����RI�C̷�a#���v����^~
)��H"
I_˃�lB6݋�%���G��ȔV��o��(�� K~N���n>CRp_�p�*�f((s��u�a�s<�ó%�˖����Y��SSx�o��S:�<�8ø,!\o��������x��[�׋��;A�2�Q8m�����	�:r+r��f�t�,m��:�Qn����@��Pj�͍�_m�N��`o���@�Zj��j3�":Y�e�/(�����`VV�'�;{=\�A)���FS�)�Ϊt���M�Rzԛ������l@�H���x��M�ϱ��I��~T�'D���2"�ÝV��G�#�Ϭ�۠����Մ/����t�lsX"]|�0��љV��W�x(�_DI�¶���l
u�7U{���$v1Ҁt�:�WF+B��@�~�`�!
�.|��QK㩔�	A556��H~�E_�XѮ�V����7���G�>�O�DʱJ��^���G��O��2�@��rM���ߘWC��Wd�N�/�$8*Zo׃��eT�Fڭ�o�,\c�n��z̽|֧ô�]���m��P���C��ej�v�I�6J򸇜A�vE�^ֶSy�E�	�Uo̉�VlU����G���������������K������Zkɏ�ӫ|�-��^�xj�H�;�5
�~�2����O�)I�����w�_/��6h�^i�ƙY��U��CW�ڀ(�/A^�i��Y�v����YS�B�:�ˇ���m1�)���Y�+r�W�_�;[�zw�cf#Y�[���M�e�BV����#m��^�S�-����%M���u�83yfRCup��s�����;�G ��X�w=���b��/eٞ���R��:�⾴�`s�ڬn�R�2����`\��8�N!Zֱ�f��u��$@o(�?��n�Cw%���H����I�׬q�p�K��%c�����ơ�̡�Y���;��g��SbS��;��zI��e�o>���x�n)^�à��A�WMSqj���d�k��r�Tض��9។<�����7�z&��j�k��ZS6���LA*뀴Ȧ�8����4��ݝЬas��#;Y)�BJ��9�GKɼ�ߩ*j%j�'߆��}��*��!l�IĲ��z�� ^�*Q(B�^�!����g�S�<N��X��U<�R����,�C�;m5?�)b�[o���^g٧bs��v�J:�ǌ����8���i1��T����jڃ�L�R�E�"��+�t gM�(Gl�qY�!mٷ�Vh���N�K�}��4����瑇�9�AP���\_�R<��=�@|lǕ|�O�݃]� 4�6��:<���}M��\���"n�b��	�~��A4#��)Ҏ>�"c�}����9 `	V����`i-<XN�T�Y�m�Va����Pb�y,��Bo�#R�Ț�C�^�X{�Cu&B#�i	Kl�G=Ho�B��U�A��T�z���ֆW�]��شM�ɦ�����\~��l� �my�?Z��v��<EЭ@�M��.�2"znq_��65�Z�ϰ�?Gm��(k;[&Y]\��C�2��V���l�	;z�Ϯy�=X�ԉ�vΕ��2������3f\Os��lz#lEK_Z�S�����~�
�c�1��q�6r�m�H�Wn����/��iy�`�����2�Z�$�V{�5�H��%�hc�$�u�ߏOj�F��f?����_��6ôQ�0L&���#K�" +���ΖL�ղ��ے�4�
��`�Ӿ	�����Me�^s�Ÿ�C�%R˨�Wr���$U}�!�&�.1����C�'�)��f��"g��fِ��n�^�̾��--V0�^�*s^���V�~��	C\�ӵ���et�w�(��4��2�uQ��e�Z�M]���q�
�4Q��Ŧb44+�158����d�W�M�K�GcՒ���Έ*G��4�{��@�gU�v/I���I��P�39���L&�!4�@��^�Hܵ�5���&��@�ͮ�%S�.� 7%�w��]^2	�/!�d����f�V�r��	�2F ]a�&;����e�-b�'��)����$�����&��oւ���T�Gu�
�/�q����5��z�[179�ss9{���U���s�f�u��i�E���a!'��W�HV�c�18�|� %q�?a^N���M����K�o�(8Ⱦ����q��{��oy-�����,�y�,��s�1tAT�yR	�����t���ا��ȭ���p�Gc=�F���A�6�Y�A��aRq~�nt~�N�àtoG��#S������`����Al��[��\^w�=��t���Q�|��.�<3!�� ��i���=�H�� ;��=]��S���l ����>����TЮ�K�d��d�I,q��t��rI�gGA��\4M��V�����g�~���^p�i#����z��!���4_�M9��DekUx���.n����8����,)�п~�W����:��|:��\$\_�[v4(/~����U�ҟ���p5�(^Ǐ9�>���d͡2]
�i*�q�im,������������>��ԟ�[^��wh�)�y؍w�7�_����rB�/���k�hW�Wm�.(z�j��?+�Ɓ���w�8]�]�t��NS�lK8�z�	7�J�ι���>�ߧOk�X	��٠�v� c{=0	c��cl>��!lc=^�����)�_\�Ӽ�<�YM�>�m7?4��6[���7�:�U N��S�x��־'�5{���l}�b�w�R�~+S���	xB��:� �xh�dR����u|�I2S����P�s5
��J�h3���������A�s��l|��/�1K>�Ӱ��5��;� q'}Ѣ!>'}��i���ь�=a����~�M�F�Ţ���E� ��B�inǎ�yM�G�Z�LV�,]IL�6$�s܏�� �p�l�x���7�:a���\�N��zj�C�u�E�rS��:���f��V���'�����
��"Z���3m�o��Y^�_n^3H����L��P���$�8鎀8�A��8i�j�MN�p_:\�7���j�08�P~�lL1���S����k���|Ȳ��|va/V2�!�>Hzκ4��Kvk�eWE�uؤ-^7z �V 90�4�#�|�f͌���W����`� X�=8�Q�"+%/��\�أ�t�PPp�D( k�3LSE�.'[D��gP�rb�p�2��Gz��X�l�卑f'>��ޙ̄a�/A�(����4������8��<fꋂ��aR������{�9��:�;�:���U�����B�-Pee�����(�hr���JCn*�kTLM�j�I-��z�u�oȚ�&#��{^ݼ��I�ןE^bΑ	�hZ��&�S��-�L*�"Q�;��=�On�:�-�e���U6A��M�k l�9�q�F�h���P+}���N6e_�1�4�$x<�+͗��KYC3��t%/>�ym.�T��5R�v)[� ��m	G �-~_�`���"���>�i���wTK+VJy�1�L�f����n.�)�4�#	�+(=͘��Lݢ��44z��U����)t�(x��6��-F�����|�'��fY�����V��&��2��zս���=^�[�Z�Y�FY<؈��,`߳i����>��������/H�kΰ�4��~/W+ۑ���^^����j����(c�o�.L_CʣQ;�	� 4�����׷P*���)g�@�%&���p.��
X�g!�	
L�w����땗��?��	H�/2n_���%%0�FP��<v]V���⊱VoQ���|�@y�j�Z<�P;`��	��d��#��h�~2{1�Z ��]�D������9E�g�4ݨ������Hl��IcA��&p��2i�G�� ����"�� ���0���qt�o������=Z}ab#'� 4_7�Z,N�&�qS;��q�,R'%��~�()��X�u/{չ�p�DF(Bn���TE��������?�lh��˜/o7S��v����xR���-����iד�Y�E��0�{������_o�
X�/�_�x�3���ͯ��g�BO��^þc>�WW�D;L���R�*�p4Ԇ\���5[�XͰ��o([ؔ�>�-&e�:k���i��JF"���e!+�O6��+�hw�n��yo�J=|��wn��`[�bݞ�;ʝ�����q��a�B�p��v����c���{r��ռG��[ߊ V�&�� �eS��tJ�W�ߢ#��H���ze2¤�f0����H���������on
d?'��9@�ӷ�f1�q˹�p��0�A?c�)��/'k�*�'R��!���/'Z��gu�*�mٗ�|mul~����p�b7'߄���E�poMV�*	���7}�G
仆���'��7��0Y���bO�H)�M{�$�H� �xK���G�o85�b��(��8ӗ�������N�*)'�z%O�W�j��\
�(@�ݧ��=�;�݃!)~�@�CH*ɥ�V��8�����Q��\S������s�)sS��X��_�C���>�}�dy��n�E�1uԵT[���o�|����4ib��q�o܋��dUƭss�I,���? ���$��໨��[�汅W��w�!N�B�o�p�XP	)jgħJ��Z����sH>�;��3(lDG�n_�(�z˯w��d���y����,�������jpŠ�~�A��19��?�<9р8�嬨[/S�pO��)z�YCWk?�l�4LP�����&�ɒ\�ͳ�H/H��-p��dP��DL�߫)J`CGw�ú�!�H���&(��(�J@Ld����FA��6|��
5𤍎�ᬲ�uA�W��=v]"�?}���&�7tC�-h,(��b��:�D4Of%��*e�izԵđ*���km�^P_�K���C�ɋ�%>��<4^[*(���H�µ�|�� �ˍO��O�MT5�K}��Q�˱�O���D��4�bLC+k�$v�li�ǌ`��VY1�����S�qy!�Iٍ��)nn��*=�E�� uНv�6�t��ܧKCX:,X6K�Bk,�3�z̾���<����"M�/���)����-
�����Ҵz����{��a�xȇpO�����_�rd�e�a�Δ��xKJ*�~4D���g�_���R�fR�7��=�w��4է3 R��� ���xE���� Y书,�j�11NN�����n,�X��0I�,�X
�| ��N%.RՊ;����M]���R�J�k�7 ��t���3ꨳ��Q;�Ƞ���z��C�k�x"����
���E	�7C�;��5s�=^t�1�����ԾXZz�ʃ2�=T��A��}6v���d#DDS{8�� 6s�z�P��Q�(�k~�7�Fdccخӱ���5}5ٺ�\��Il��'=��	�DU�P�b�*a�KhΎ����	.G��u�&-5���:��'�-����6	� �Q���P��Ư)�`�,�|�},U��Z7b-tQ`_eV*����I,Z�kA-��-�89 �q�3�&�F�ଂx��c_+V[l�3$�ulO.�)e0�!�~棹�Ǌ�Q���������5�o4�dp�oFH����R�;������u���L �	D3�K���]���^2����^뤫�0��B�[M��j�_"ȸF��fX ����b���r�0�۲G�+n�ښ�t���n�Z`na����k���<�����U�����uFy�� Ym,V��Xt�Fzݙ��z)h��*5��#�(٩?޵so��y��&�C�"�#j�IΊ�/�K>���� ��¢�|.��\�aGZe�p�ݰ_0ӓF���{x6pi|؞�ْ����C@%Az��/_���Ҷ��[[�gZZ?4v�<R�*��N�s|̂x�2c�W�53BHy;m��<���Q�C!�$!`�Н���l
��R?b�p��G���^*�2��kw	TF0D8\ET��g*oR��s:��\R߈�V�v��VTɅh�hp5���2tZ�D�n�l���������Ҧz�wS���^�81��pB���	��7�K�kJS�2�joV<��W�{߿e��{�d֖G�R��WHH�-)�,���>���Y��/]H#��
��%	�Q+�`�Zˋ�6��mf^ˢ��H�;nϸ�.�rC������z�U�>X�7+l���g��|W[ZcW_���GY����t���V��Ӱ��w[(f���0�E������
�=��+�Z����]�_�X�:�Ց$}9�O"T���$.�ڦ{� Bn7�I����.Ђv~�X�Bu9�/�ȕ�������B!_�k$y�p�eq6f��e�xJ�Hg�f>l�=�@��r㈂��<R J`|?c�4����w`�������� ���S�9��İ�=��F���Iߔ�*�dMaVX�,�_
*�o�,ˮ�o.��*�5ƫo��"/�����a[�s��0�+ݔ���ٕit�k�>:�r߿���]\�YV@e���⧣Ib����R>�q�~��xLx����Ж�T���Á�}�J�~Mښ�4=��ʬBn�+���fR!��z�z]��3�Glƕ.�gY|�yF��v]����s�;��rm�< �%�Xo�W�B�!�M��qz�k�lz:� �N��*9ȟ�G�$4ZA����n�L�	�9�#g5��dIo�	��_��lE�<��c��ST���@�K2�`p�����C<TA�+mڳn�>r�@��ȫɮ�H5�������^%[��*f@��7iE
��f/MAfMȉ �6M�R{�f.Ú<B�\O|
�G�!��%l�H��@E�[x���`����1�]�HӲ�WS ����i[�gvZ!7k���TB��dԓG�g����d�s_���~�Dd�+�x��%�Y�Mr3��M��~,��`,�,��][�=9a�#�.��><�w�-kؖ&,T�f�Z��
�_���59�F)����P�g:�����hFq7au��z��>-KasN��>�����O��F
�|��2���
9|&��<.)HF:�nO(W��w��$r�w��FS���oJ6}��`W��p���٬D�5����J�	�X�����b]��L���d���*�Q�b��� �'��0�:�{ atg��K���X�A1쾄r=#�-���p�X(�	����$y �W��e��ArJQ�$��J-���3X��������me޸�|����f1zJ��ZG�%�>�;�]d��싺�Ҿ9��j�r<͠���P��R��[�)�6\{�K��;�t���
�k�bү_�z�(�� Y�*�u�}�H��������~�U�|v�w`E�G��ap�vڛ�o��z�"m�g!~�V��T�7��K�۹1O2��a���F���dF�������q�S��7�)���J�Z�eu_|Z
�f,������gV�y����",�G��p���A��? ��_(Yz��ù��,���M|����"��:Y'_˺�ٲ�	�M�wb�zO��ZPO���0�?sKj��1FⰭpw�5�����:@�I��d����j��r,�(����M���}B�e-��{ED�O4�?��� ��Q~ţ{a)bU�-	�aG���Ay&��ZK�f���s����߾��'���AWd�'�+�����_'�>%;І�I!
��'AA\M��5l֛�^�:R��0�@��x�*�GY��®��$�k�J-�}�[�NC,e����.���8�5��֎���ڹ�K�l���Ş/¨�8$�����ů��M��׀���T��C2�cp?����� � �0?Ì����:��aì$��2���9���y~Q�a��t��[9��E�$�7f�*�W�l�;j��Ey� ��E�"�/��s�]�_f�G�"/��!�.dR0�Ax*�B#�$��p]TO��OVJlB�h����l����>Qp\,u�S�	���%��H�dm�7�+N�G�,�D�R!Q�@��hxR��>��w4�Ј�TY��#0��ߌNk���x3���U1�YE,Q���&fu �=�K~m�гAr
�z+��1��J��Q��Y!8�i2?�U"��ƞsA"��d�N �v��#���v��e5�sKH:xiJ��eg%�O��ĕ^1*��2��B���>@rq�ڄR4�� �oP���b�y���3?3��'Ej�]W�Z����wK���]�b���B�jl�7�N�C��Kh���EU�����7d�f?��5zF2�xX���-�B�ʏ8������5�˄����t�5��K��=��odlȈ�l�w3���p즳P�L���T~����@������:U�_w�7��7�n����'q����L0T�/�~a��(�:?�b����>�S�^n����O��%�^�T��s��������Xd�p�|U�E�R*�	\�t���;��7&�cWd+����r���a:��O�J��%��M]RV���\��*��}�ʙ�kS�6�S+t'��1tn��q$y"���C�kɣpjm$�ƾ�1��s�Ʉ)� I�>  ������%c���,]*�)`2z��j�͚pn�~���l�~�`�#�7I���*jY� [��A�/�h�F��] .l�$/�2II�B5��a�4-�?�x�8>I�gYc�Rjy�&�ڥ�7��ե�'���'�I���[D�Q9��-����T�4����#�,�ߩ;dne�����2v�J���`:}�t��N(	�Q&:��|ܛ��L��D� �l	YY-cߟl�����b�ҋ����L%?���-Fq�	��3၀��ꈖ68�΋S�<!־0:]-�jn��0VŁ��b��&��ȶ�!�	�i+����/��m|<�f?$adczXY�����Uv ���$��mCW�<�v���\;�
��f�%b���7�j޲���U�7�yK_e^���pކ�a'��>1�M��fu�J�{�l �(�yE�KQ�5u�Q���Ƣ�-N9lz���:=� v�>�^_��1|;���E��$�(�:�0�`ٜ�`z�Sy�F�3��p0�d�%͒c1ȹ�I��+$��o�t�=d��hE��*�q��8~e���7.�R��G���q��,$C��\+��В>�B���>#O^}\q��rO�`��*����
�Mn^D�쏆o�q���^�mb_I���`ߚ-p���U�&���O>����ӷ�^��/�+�iڹ���D�����@�L�"9���i1�����}��>��C��r~�t��?�L+=E�HÐ�T�6�<�����-G���Tf��bX�|��7T��_�k���1� |6��r&Q�\q��������|ٴ̓ �f:�3J�)���V���DU��Y85Џfc�<)�=as��<S�z�웝��_g:�Fi'��{)Ұ�;�>N�R����I)�������#JU��:��,�Սr��#�J��5-OW�o���B�:̃��Ib��[c�b�bB�\n6!+e}�e�C.�!�_l�B2�Ra�)���P��jQ�\⇟�J7��)1>����f����`Eʣ����hLAbk�ύuM�y|u4kh��VR�q�v��gZM�]|�0!�Y��Y����-��k$��ÄY28(3�2|��&ΆY΁�#������<y*�X]���Fj��Wo@,��t��w���#kiՙ	Y�+<j��t"��1�V@�p�F�x�6^w����i /8i��I�5u~E*�I����0��D*9:�j�K�(�ތ5M��Q��������s�Kb�����36�y�>��7�v	�BJ�B��z���� k�����[g�?..��� B��%�@m��{cZR�Q�٧Y�2EB�_[]/��o�k-�.#�U������p�5w���-����}nu(���$Rx�����z�@�E�Ќ�t
5�<T�/�A����yTSq�A/�h!փ�����3ސ��d� �$�*U�f-+��j0lG��S�/U���tƕa��6�C1ä��7ٽ�m��H���!�N�~{#�_r�0�4wA�n'�<u.��t+�*,�4��af�8Ө�$&��*u�(JƍX
G�C[�n���N2�og���اh4f%��E���2�S��D�O�?�+|1P(�)��J
e!��.�q���M���Eg����L*4�b���mOϽ�Ъ����h�}��[��aU,�_���Z|��t�2��~n�⭏����WT�h�ʤ�	i�7 *B��&) ��ϴ��b�7����S���f)CUT�����nK\��]�G�!=8z�����MV��Cݐ�ϣP�7
Ꜩ��\��1�_��>��
��p��|/��A�1�@���_��GiP|oiMtV��@��+�Mjf:3z\���{�O;f��o�p�U&�$F|	�A#���_;�A��"��:[R|J�e��pD<oV�+q=`�p���R��E�W5����el���׹��c��3�͢���`f�R������b�n�Ȝ�� ���,���qtk|���>|�+e�d�ys�!$)⢧��3ꡦx��UEa	��2�~.d#,T���^/�,�t�o�
_��-�Is[�	� �s"E|�G�(;�I�]'��%+7~����5��s�2'�l]�!
���KD��>�P���bW�Ѧ8���	��=�mi��X��Dl~풥y�����0�X=��9TB�DVT�6��&;VfVF�)%>�l1�H�I�j�"�ԉ�n���⧚����!�ݜ:sB���?���e�3|��GlW�h�'�L����5{;=4��×�����Ԍ�җ^/�u�v�E�(&���N��׸����zBF���]�B�9̈́��^�z��s�J��\��!�e� ���u�����3��U�#���r�����m�=%��"d��(�l*��%����%�����X�Y�?ӯ�M���7�U>^'!	
�����{���7X̮�~���"�⏕ϚtI�+��&�e��'�R|WD­�i�vwƽ(4_�f�$7L�տ�h��1%�۰G�(&W�쵣� �}��U�Rft�$���' �b����%m�u�$-�i�������pfV�Y�f�]}hU[�����Dw�u�ʿ���B6��*fN�8K+X��@�{��ra��D[�l��0���Wz�L8X��t����#�&J�2FϏ=���}L��ꐿ��{6�-?+�+�j_�z�E��?���:��!�í�X+��+���3L�?4�0l��K�!��Pj_�Q�>��~�;�F,㝥ȣ�������I״ A�;���0���Q�I>��{+�${^�<��[�ɋ	��̓=��n�2|�����/7�Z��
�	oAaa�a�N7�p���j����S�qc�y����>
"�0,�Q�Ȕ2j�9����Ӛ1-B�-�P���I��ρ�͘���`< �����*����ǩ��OI��H�� Y��m`�ºb\�!0��Ϧi�������\E��D}<9��a�袻_w�̧Y��ڬ�~d0b���b�e��ijB�ݗ�D�� +iWD��֋�T����e�%(-��������5��L�/�+��F?`~f�[�!�LOZ(�s6�O��Lq;��ȓa$-�?&s��o "�䆩�q���T{h��m�`�0�4	�c�=���z�|�F	���՗7%0s�'J�uQIh>���QO@� �3.��}��.���w��+�	 b����%B;���-�3�rr���Y�U��X�XIv[�0���3�odɿ�Afzy�i��Ahg�)Aa-'v^����յd����=mI��*e4z����s[{��k��@B�rW���o�Lz65���7t��:��\O���>p���1�2hy5���#^�`)�y>1y��n�%�.{��>c"72wW-k#g�$�e)�0#p}��5��ǥ7Ś�����#!v��a��k܂P�7�WD!����QC(a9nx���CɃ�YƋ"����&r��.e֘�ѽ� +J�B�}!�f�p3��4-G�0	0�Y�(���~��_m�36�
��N�����g��^�z��I�n�.�Y�_���$�A-^y������O�7�Oq_v��U�ɾ2G� ���sȂsb�C<{�\��5�I8N��=�Os��#����b� �."-JЯ,�H/A�4�G6�B�v>�SZ���g��Fm0ok��[ì�s}vz�bc����ȩ���a`�}�7j�����k򭀲S���A�1�[q��_��ŭ�7�M�)�Es�dx^^G���Ac�~WX�˨-v��@�Ǔ�6](��A�@��y{.|�-��Exo�:]����+xS���v�c#@�)�Ņ�h�N���p6��%8"7��l�jnU��nr�0J��O@��6oo�DWJ���.W��O���&��&'W�h���J:�Q��f����9�(�,o���9�n�F�ʖ�;�F����o�-��|$����r�$|n�L���U��*�P?���pK�8���_&#�/t�H�K��c�f30��G#	�)�U��v����[S"6qx���=��$������D�����}��C�A�c�K��6Y�Ut;�S�ާ��Uf�b$L�I�
�熙q}���P/Emꬨ�u���/���T@c�!��{m���iW?�C|#�����a���{z&E��if ��9K����"�XN��e
U��{��XO�K���ѱ��W]J��X�	h m�ex��H��Rv��V�;[�Q��^	n���t ����d`a4�:��y��,cW?�D�	�?�;D��M���
W��G���]�"0�]�b��VT ��X��![(w�U#��.�)}�oPec�t||s>�po�"�����jS��ڧo�p$+��k������V�u�n�:��t���B��<4m�|���Bh����º��2�˖�|��~py� ]��˟�l�bn@'̄H�{=!�qSY5��.��pt]LM��p����1�=�^��2��X¢(9���D���
����O��Ҷ��+����ƕ�k���w�]A%��� �iã�Cx��TP��}v�W��A���Fh\��� y���#v!��q�?� A'2h�����Y�Ae�YT�2���='�6�c��f�3���g}JB�s��5����p#��p���R�m4Cw�
P���`k�=�ȃ(
��|g�!T���[G�"+t��wˌ}��|V
��X�97�JkE�m;f^1���E���ݧ־�]{*�6�K�z}��[m^[�!f�&E[��M@�̟+�,���@�/�VR��Y���k�����xZ��tI���m�k*>r.��=��|�E,:����pz	�W�-�z��%�r[��zԌ�I��.�,g���BaW�9#=J������/d�7��݁#�z�*�փl,��]a����gE&��XѴ�_��5����[ڗ8�7P�8�j��Q�� ����f���T^�Y) '� t��kyb<���G��r9�ac� �Z�����HWi��~�������\6���#��y����r��!�a�rk)S��3�Kr��0c�F�zL�O����Kݬ����m� IF���U�S�6G�3���p�S�!ˁr��)��}7΅���r�i��7�U�1����x�� �+#t@�U2�ꌒf��e��n*�GE��\�3GC8Q!}�[����^�3z�7�Wx�9^��0�0��$�퐕E�ry,h�w�舷V_����M$����A	>����H���y�|�D{��Gt�:�]�*<2�e�kMv'"��X���q����1��e8�
�N�����fi��X�FEs���ng��]��v��R��ݿ���u	�cL��4 ���u�9�T�7�j��I���É��=9�N����W�t��xٛ��њ����-���	�3����:�ϗk3��}�j�[ǘ�%�X-��ak���PÞ�х�t�q��5 �� dy-�A��wcicS(x�<ț�����D��`�����K��'����5�F�"�6��Y'#��C@pL�L3���2�_�װ������X(<y��h��G8zhm��	���(o��0LB�;j��\
���)e���P�=���yE%��PT�����:^Ty��坢�#xƍ�>��ȶ�>~�2h�?�ǭ�F��:�O��2� ���s��生#��1�R[ֈ�&������x�� �0��`���r��Bo�U�GhH7W)����B�۞�M,;�*�o+��$���.��y{�2�T�E�I��`�WIP���DT�s�j�0�nק(Uj�]��O��x��`s�.��mtWxά��0�4������Z��w�=���1��q�F2y>^m]gL ��p��Sź�O��/�B@������?�W<?[$J��g���D޾�(�W��QuϭO'������ްӭGfvw5�[��[˩(`s_��hF�&eb��s; ��lSچ#�mB	|��V�$�pE,�ǆ����rQ*�.��	Bry��#J���5��P��6��=.�/��lɱw)�}zb���5�½c�sHߤ��CM�(�Q�w�mJ���o�T�=�d�Qե#FZ����׃t&q.�O_�w��u9�$��t��K�� 
3�R���Th���٢�xo�vm*
�x�Z�i�5��unY��yT�PA<�����
��ű�۬z�r8��B;ū�;�2AWx���[Ja�ie�k1s�>e�Y��b�sN����N�Q�J18�ڄo�t�@���73�\md�L�7��qP��%]P�g�_i7<�'�k�ɛ'���@��l��ǆ(%�gR��X��ԅ@i2�ث��#L�$�>���n��c��b��,�I'U�b�a�3i��S����1��K���cog��]�<�s�Q;xc ��IYI�8�}W��|�F��'� ݧ�U�i�Ɖ���;7����Y0��1�)�	�Yg��h9x3����e2�����U��ک|�k�9���=�L3Vt���BRx���Dp���-�r�����S�^���}�ɽS�~���CBPt.>#�:{���mn$тt5�*$X�<����m�������z��堯��4?"����Q�L�,y=8=S��N/�3?��"k,���P)@A���d��z&�0�0���)�|��<B+�.��,nn�}#���K�
�}`�b[��r�!Y�'���EZ#��+������	��\r��څ	]�.�%?�ϒ���V������q��Vi�󌘫�/l�L�z��������R�a�Bm� q��I]r�# �۰)z3��9Oe���I!&&M�h�ᆇ�_�2+8��|�t��|I`S*�6�{������+
�S�H�ko*�p����� h�����8����)�^�������DX�lBA� �X��RZ���]���e��!�9�L���^,�S�����m�� &Ĕ�ww��#U�Pᮝ�e��<-W>�d���� `���d	n��Z4P���������<Bk7Mt9�*��Ed�!��O1�kF!�@j�ĉF�2��O5��+R��`:
ݐZѻ�Q�W ��Re���K��_�$�E��ݱ.�.�,��[|��M�bk�!A���y~yW6�� ���Y����ao��=�'�F�k-���;-�)4'�բ�=QK�L���ݤ;kP�,aբȺ�����1��<��!���F�vY�����y:�*�&��&MƢ�0�q�7R��m�v�(����Pa`v���S�z�����A�>���#��zi��br�`��Abn����F^ZOd@-����&�C��My�u��(y�kv3d�e5�u�䫎�t,�g7�?_�p7�W.rS����W�[���̻�vc�L���D���dN}�、j�
uz*
��B�?Vۃ���h��$_:O����}�t�����Y��3q��܌P(��{kY!�w{X�`��5x��G)��*EX��1XN��aR�~ʚ.��,��~C����U�|]x �+qg�h��SM��FzJ����}�^+Yd�U �1�����B9�j8����7�'���H�M���:�b��b��P{����G��3'���@��fuЂ����N	ʆK�6FuR*���\��dE8}LTc#S���qݬC����F�L�Bs�ma�ۧ���y��J�q��&��rzx&s�@���t�g�/ѳ��ˋM��e��wĮі>���S��W��4��E"�QtX�t5��x�k�Zx90~)ɂ��=��XF��b��$������
篣�S���d�a/��h�3����/�Ye0�������=��S�J虅�l�����\Y���xD� �q�a`��iS�lMG�k�"�F0��=W�5ױ-c�b%�!n�^��ڳ0��.�r� �q���ũ�t`P:�Fd�܈����Ƌ�;T��O�ai���|����l �܏蕚*aڤY����D��Ao�?�xZ�v���[� 9������@�1���	:$����SZ-d8���P�cشـ,	^
C�H	�jo��OD�a�6���f�x.��(R,l+1a���>3��aיI�f�? W��A<8C2�$u	��k�3�6lL��Ĉ}�����W��nWG���ezH)R���&���0���Z&���ͺ�J��j�q��v��O����#�>�ab�o�N)�0�}Zы�7�t^��c�1�T��zL#��%ʣ�ް	W~?*B��xGE<��>��!���_UZ�Y�����Є\�WY�?��'�.��J��\��H������YG�ն�:����{#��f���w�X**��d����T�
�u�(^tU�GD���Ĕ�.Qم��d'��d��Aj�̂�@=5�<G�W4��%ٞ)R��ٿ,/;�GB�/���Y;��)�w���r�?��٨�7ckY��5R�%���hY��W�]�D$3�#[��[�t~i�S���V!��&�?c���'�߄Shdc9@pDM����#�W��	��mS�=ƾ�wT0]�U��Da�1H�]9L��$����7�ds��/K(g��w2Jַդ��M3�DЍ�ߊ=u�`A�X7�`�x{�α_X�4;˧v<^���l��c^.N�Ȧ����V�Vi��H�(�&զۍ?�a<�A�ސC�5%����na�G��ל�=-�t{�%%�^b�#����;�v���a�t��2�b7��
J�Iat7)e��I���"���z�|$pQ�˜LuA��	�SWL|ر7�2$lBk�N1�H�ˏE\�����S0�ra�?+�=���Y�z-��(�G2�:aR8?�:B[�RQ��v��&���+��W��rSc�VjV{���N���X�M[�"����S� �7�3��iB=���Ý�珰�X��g�?���WJ�D���	�$Cn�s����񲅉|?9^G:R
k��?���е!�M[)��
d������6�e2~Q�F�G,$`ߋ_N���(��݁c�_
-~>�\�ڀ���oP!i/0�ˊ��ptV�s9V��}h2Di�/�2w�c�^¾�L����b�|���sP���zq�˹���D_h��ౌm+V�N�ۉ��$e�%m�C�`j��v��� ����'(�����bpC�\�t����|S
,�@�Xu��q\f}L?z�N5G��2�wJ������C0��/��o�D*%��k�dG����g��Ϫ_Y��nզ������`Q�P�>�G)��u32La
�X�H�K��I�TVU�����þ�֔���sQ̵�q����R�+#����&���`��j����Z�/������S�_�w>l����%����2�%���A�S��]�PY\[�TFjb������������=tߞN�i���M�����a[���6�FS	�~{*�@�"x��u������1g
O���ʸ��[<���r��O�oSzt5<U|��4�b4ԗ�˿�d�zd�t��.NC?���}?�O��=��nHg�c�>%hg��;ܿbZ���s_w��MUMz������eRp�]C�Ƽ�\��:���kd��効����ɂ��
�lQ�꿙w����d�ӎ>W/l0�7��[R����JB�p�fh�{�/��>�T�,�D�G|/���6a��v�b�F�\�6ܷ�q�o�n�S��:Z��$�-4�$�Y�R��pނ�[�#:�,bH�Ac)�@���+��CqZ�JN�����-܌��;�'ڊ�7��B�[x���A���+sS�6�^g9�ɴ�C�"~D���s
Ɂ�$�K<� �F���So����Z�z�Ԑ�?J������S���8��X���Lj��Z�Q��&Y>�W��)�{��*���r��0���u֫T�$SVeT�.J�w����_�$�.}��b�l�]:n�J��ƀ���%zR+�Va����1-?}���+)���s��|�j��`Z�y�*�BZ�_pZL�����j��F��������@	�Ůe����$�̣�/ ��P�b`�R#�X��[P�Ҧ��0���$@1���[䁇^�b��8m��'8��z��G�f&`��x�Μ���ژ��.7i)�����=N<2Va,��?����{�����|��A�Q�T���������m���G��c:�:��*��T- ��ѡ���������a�$ҩ�v��:�]��yx�~�j�st��9 �VBNO3"���l�d:��%#���/�h[;Δ��-� 0t_l-�v՘,w.d��{��ã����˭�<�W;�UΫ@�.�g�@�s�<������u)a���HB����(x2`m��5���t�,�(�-b�㉋�?Hl*���
�_9UZNn��O�D�T���^�-��kb"E��"�hJi������e��3$�.84�n ��O�c��/�<�$����'��ş΄� ����G���T�|]��bYI��+0��M��fj�X�����?���@���U�Ga�˨�)�Ii�p�\t��0�GÕ���p`{���V��u�n ue������V�,1��"rKXVR��[���M]���r@�MX)�'=����� l:�>��M+�1�4��8�J,V�L'F_����F�N��G�'}�C�P�����Bգ�W����[]je &�E�=�#�t��3����23{������L�V���&ǣ�j���ɴ37�n쏤L���&��zv�mǁ	�ߝ�}��zĦ?�E�Mz�=4+d��)*z����}h�m���"h^5x�Zb�FrS�'���ǔy�m�ʈTR`7<_�]<��Rc���M̧|�=���0�y1�5�"��_�]���Eʷa.7�s�#"6��+���A������˸��P��,���#�F$B,����)-L�f6f>m'#'��a}ְ�]��� $��T@���5�Q���z���"�q�)�s��('�Z���c�1U��6S��q���EH�(o�w�F��{��#�E2�9D���-7�Tiݣ�Tp���t�2�}k+��V ⫬S2�l]��"�#��1-ܾL��zu$J��0�:����F�#��@���5T��*�&�X枳�>N��῜+�E���A��9Bc׳��[� ��W_���s_v`�xՔ�7%No�M��;.e@T-���$	J�|��l.͛G��f��E`�p���2�/�(���2L10M��vKh�"��9��"���;s����@���;�����*>����� �����oϼ���T�dG���s�}���c�TT��)	�2��eM���j���b��R;Ivw¤�C;N拟��y�����t<��Gӻ��u m���)�8+�!���-S�1��:��ڪ�L�WѨ�=��K�H�	t��@���VPk9�I���n�v���
�6��=��&�g�""�L�#��u�qՉ����Jw�:c�p�/�d�ңs���_8�� �Q�����ԛ���B�M� ���9zv�`\�m��n �{E�{԰��D�nk:v;�ܟQ��O���0�,n�p�����R���z�Q��r��h> ��$}=���h>�J����)��1Ūh������b�l�M{KXFP�}'f��Xŉg�Ѿ��
�Y��y��Yb��Un>����F����������֬`�cf�e-�p�!z�W �4(���n�h�,��%С�ߖ�v���_�[1
����s�Ỹ[��B�.8�4(���nV��B�Uo@����Q��b�T*��1�h�>+�Gl�����N=��-�	9��0Í/��ϒ����Ǵ	�b�1��' �7Y�-��N胨PdC  ��쏪�}	���Y�8�B�m{��z;���5�/�E᳸\z��K�����^O(�H��u�Q)�k���n�ڌ� ��3s2�J�x%;��E��XO��x����7��ˀȎ����֍������"����#���b	�/���`/�qK i#�%�A��D��;>|�m��rY�[�C�K8�g��RL����/�¾Ow�뷊��䑊��E�p�|#�_���~��A�_�2��tVO����H��Mܧ�/��u	��;q�+5�������+��]��K�Q�Y��w7뗑$h5n��`!�Ik	8&�yC	P��xZ���R�� ls�*���^)f^IH/*���l�\ٞ�r�x=8w��K�UdwQB��O,1��lB�mç��/���4#!0�JґL���N-=S�zQ߹���p�q8�ɏ���I��(#�%��y&s]�`#����:�ĸ���k���#ڞn���Q��:�Q�o4�;�j��sl�xu��癩�JȨ�����6v��'�3��-F��i��� F!Y	����Ё�+uB:h/��mJ���k6�����V���S�:ut��L�0���r���}��l�̬ā<#�l#]B%!��}qe��I?��F���Q��p1�:��������UZm@�w,�5�E���N��E�����
��&��яh؆/�>�.�k��䘵�a �ajk`�U���o��-�?��N�$����Ki���U��� ukF�T�	߈�AxrYM��������W?	���������i�`�o��|��~��̲���,��@یB�Uk-��D�?��>���HB�})sF�Jo�o�.�|���N��PT���c;��n\�L�.� ̷�?��%���W�r5��X����8��_ǻ�g�`�#K��*z�}��׎_]r5o̮�z��IN@�;���0J�?S5�c,|�$}��z�Q=Z�rc�"~�!*h\���(��9��kbD��ڼ�fBOw� �+�H��mMM�!ht���A���x����G�p���N^�7��}�d݋O@A�T	�.(& �V��#�}������e���Ld��#��'�" 0����?�R�N��6:I�匐>�g�<E� @O����P����5ԯq�_�Y� ��o�Rs���#��L<�v����8�H���K,�Km���|�� ͑��7r��
I>s��$
��K�0��u�L�����~&Y�wTA���"�E�H�~��{�՚�`%5܂���̐�l�B�8f��q�$,���l� r&$J�t�f�N_��7��8;K&@2w]aF%q���Xw��HW�U��'��?h�λ�;�Վj��y M��(~1M�]}�/�B��%=N�K�A����^�Bh�X��J��O{��l1�k�kr8%H��8�Wr��&��rDW��a�6W	b^��j3���]>����]�I<��6߹&]1�ᾀ�a���ɂ[J4����(�!S�%���@I�JI���+[�ߔGD 1�������j|����E�G�-�<d���z�Y\IsU���9��X���z��c4�m�ry�ȗ�V#}���1�����F�j�#�ۤؖ�N�ڌ����jx��omJ)���_-I�� ��t�`�G3�y*�6�z
�YM�.�`MP�l��侢gF��\����@����h,�|�F�#5C��D�b!F����� ^���o�̈́�d�ö��8(R����.�J��&���$�Q�,(�OXR�Ў�&>z��EF�W�scT�-��oFۼV~=p�K�����;t�V����8���������L�UP?�>[�-���Y�� k�����ϪHF*>6���n4��x��@2���w���C�v���?ca[��U����7Ы2�����@Μ��06@:o����ƻLY8f��́�i4�([�h�fU��i�Z��,�s�7qb���|�.i
8���e��P�r�Y1yXW�6��R���y���}]��r����]^�?���j���3�+�������Ġ�v^���j#<|1<��^�	Ѝ��"b�.��M���.�[�S;O������7s�W����O�%T���Jv/ s�oe��ƀdU�||�����+X^�jҨθQS-IJB%S��Q(q�s]2b$_2���TX������'Ͻ�2�9U6�������l8�f���rH~
4(�2�����:h���Y�1��CG�ͻ�f���%��v������~ggZ������!�n@Y��F�(u���JnvhTN�Wp`��LX�Ɉ�p���*�x�@���xRvm�� ��������׺�VE�?���Z>�1Qi�Xfyt�!/�!���g_�FQ _�s������U.��bOH�w��~u�{ED�op�;�a�����_"�������(��x�n`)2�wxn7�n)�$��_�h(pyu���؃�"�"7ɿ���2e�ɏyd�\r;4Dü����fK�.���a�����"�sӾk�>�l����^9"�����L����'([T2��bE[�����];��DUQ@X��oߒ�Ф������Ι�
%R����w�$����`qI�JÌv�=?qa6W쪓��<���4�_qDQ��qf�du��?RQkyX��=�+6��P��'����[dɕ�&���O�v������­��@`P\�b��5F�y_��6�a��
a% W̍��f��-�x�B���M�&�}ڪ��ꤺ���l�,(��x�6e9�\vsU�{���`QTf؝���+�}B�ϻ�."��o�&gڤN0+7J����e�s�9�X9��'ƚ��:@��j`(��<=dk6��̗h�Rb����ZVH�24\�d3C�n�'!�k��pB��ȯm,4�9��0=ofsi�ڢ
��;��>�kx2����C�?�.�� ��?��M�����;-���q7ylnO�U��Ww��0fM�"/C��E�D�Qu����B�1Y�^�2��+q���~�*b,V�IĮ����4p���t��go�r]�ݒ 0u�+��D�J.��Z�mƨ��3�T5�O��O�-�d�~�xZH�q�t�?AFa}h̐��0[IT[�����5��2�de�~Ҡ��i��PE�v�M=+�L��+�!֫��
Z���H4pc3�k�����DJ!�P��M;�*�$�\�g�r��������ƅ�jT��MF\S=�|{I�'m��� !�8XQw0ɠ1G���,�+A�������c�"����\�n�S��� �r�|#y�q��>.�j��A}i�O���4�-\y`���/d����w���2^�OƼ�A�N��:]-k�b�?��F��㏹�����W�̥���!�	��ug����oZH����ĉ�#�9�[�Z�����j&�^�Wxk��3�3gr�>Q~�C��4%�7�Ғ���R�����O�Η�(�e�/ț>��WBz��r;M-�G�ۃ��:�%C�r�^!��ct���ME��vdaz������/��\9z<Ak�#��J���W��4H[���2d�ji��=�u0S���Y�)#��5��|Q�+��ׁ�^��I��X�o<��s�J�l47gRQ�!C���!�sq6��2�5x~p97$���hun�oh$�_d jR�#/��Ħ�D�%sX˝9�i�T�ߌQ~m^\M�`<D�e9`:��Qy2ㄎ�-U�#ޭ-�N��C�<^�H7�l���$�9��W6#�����<!*��I��k� LӁvX�I!k��������U�^��*�[����/ ��S���W�B�LZ��l�����L=��~�#U� $K�X(フ������Y��BiZ�i����pZ�3��2Z w=��+�m��,E��Z�m�����Sy���Ɋ%���U�or�![d��T��K�׍J��{���Dϖ̝uz�DX�[1���I~�F1�3$��|�Y���@wA��[y7F�7�SD�l�H>����$RB��6.@��_���e^�4�\����"��Y�>SmڴKb��1t�u�l�)�K�\���j�@����ίУ��j\`�ȟnЏ��+{ųl��n�/4ZN��?��!i
G�I"qU�@��*�{=����ɳ-�s��ה��99�7?na&���P��B�}#��5 ����r�*E��e�: �����Y��2Q�2��q-��5$t����B{�]�sd��C��pr��SCkb��E�[��B��Y�vu�jP�:�����D؀�\l�;�5	C��=��&��,l�1&6:��L�(�C���p���g�����#�	��~�3)����XKC�jR7�B_]��x�3M0 [��O.�)2k�J���H�/�oUg�W��p�>�s�5 X_��Ƈ��w]&�EPEIp���{ˣ�Mu�f�OJ̈́��p�_�".�}���>ŷj�mRS~Rb��fjz
$�/��R�م.=��&v�*1ϡ���C˗�.Z��؂�p�Է8�b��e�����v�o���N6I�Kܷ0j�:
Vtz�U�j�ٟ�r}�:q#cB���MP؁U��K����Ǿ)۟px;�>x��iY��2S.�/"c�b��\���d�Z�^?CL��R�(-g��]�o.gJxb��>�h�3�������OW�u�)/�N]!�K��5����q8'1��aB�v'��IP�
c6��fD����[��BG)�w,jҵk���oK���IGs��ͩÁ�x�銱�RZQ5�i���L�V�Ơ�5��cS��0b�O�7�@fK��ع����������i4K$�5�-�[ضB���,��,x�;ܞ�~�����m�8�E��t9��?���>b��<vq��^�?�	��>���vUZy��E��,�!��H���/��O���nʧ�ِ.�Y9N��zV�Gy�]Z��wI�T��jy�;_��'+8�Z7��X�Z{�Jϛ�
�����R*�-LF��$J�kmn�Pş����_ğ�d���1�6	!��o��3�(���\��/�]6Oa�) -*�}���[X�<�#vB��"|:nل���L�L�)W������)^E5"��q=�����S0avs�4L�-�u���JJD�S�+-���7��e�1O��ɑ��F��}�<�!�R�촃�;�Z����:�a�I�6��͡�/]�}�mk�,���5�%&�e�&(���E.�����%
 5��������Hc}y��]��.������nq�m�l���i4�)�C�����R�TQ4��P��&Q�z�*0d���]�L6��m�nm�$�4��Y�ﾍ�S����$iW,}E;w\��6|�I�X��G�O~e�� �������8o��qi�'L Ѐ[�s>�6��i���[Ί{���ٟ�Y����.�Z�����'�k�����VU'�tG78L�+�㼁)vqtC��uց�W��X){)e!J�&9��ގ�Hc$�� 'C��@��*8u�3=pЬ�/!��"�� V
��O �҄�t�X�ŧ�b���_������ ��@č྇�]���gΆ�5?j��G{O��V��?o���a�Dq+73D<3��3�1CHe8ݷ��Aгˠ�o$�\���2�Y��~W-^}�A��u��T�(�?����ũ�3F�Ň����Ȓ�W�虉1_�f��߮�y��v.�ax�_ƨ���p��-��Kc}I"A��^$*W8�3r��1��)c�㎖Z���3pՕ��`^�=N^ia2Qi��o<����G��rf������7���Y����p"��}c��|�?�:x^�L���3�E�����y�$x|o�|E����D��}�`v�bs�d�`M󫪟�������s�R��h�@׎<_G���Db=$���Rez��H '�`�D��$�~�kg���k:��|� {i�$���W:�ga�7� 0l�z���DH�e�3�딉U!���ʴ�	��X�5����Gp��Ƣ�c���'3��
}#^wj��K(����n7��5wku�+�R�ϵ�z�H5Ô�S�U�d��ւ1t�m���""ߠh����"�mb�,�cf� Zqg�@E[�I l2³z��8!t跟�o/��/��T��Nh�)!��k���/A��;ͮu��ɸ�+ͳz(�������쫪޷�nշo��T�������j�
�YX�݀�M�ù��ʔ�����u�D�)�^�<��X�v_)+�ܴ�V@�_�W>\�4��o25�y�
|���i�2��,u�T��pj�:d����o-R�3�� N���y ���#�d*��4���ٺF=��=�v��P\+& ~���0= ��9�Om�ۤ��v6�a�H��[:��n�ḑ��k��MHK��-�����Jf���)�����T;�.rG�вEO��W�S���� 0��P����ѻy�X��0#Ⱦ�>���ˊ� �Ƀ!�䁑K��-@~%�g�O>�[8f���F �*Jc�^���I�/��ˢo�#~0�0���MO�
2>�y`���Jp�4�X�r��$�҈m��dY��`��Na�W�����B�Y�l�9��]�G�e-��h?����He������(�p��Px���5gp=����::n���$��=ݛ�-�t���mѴ�`�e��*�)Q.�D���_p�8�3*�o\��ۋ��]��ʁk�y9��ӎq�[w
�H�[��AD�� ��N�/��ɸ����/F��nOQ����30�)���Mڪ��E��W,FP�M�~�u�c�7�_������AO����&[}�s��@��^^d�?)+=��55�4N�c0��%h�G�߇z�tY`�G�^w��t/=�X�z�)R�J�7��W�?d�5��|�QLn���x�M=�J���3�!��{TDC���JlҢ�A���:��`+Gj~�\�������*8�::	#�<�C�g�Iv��c�]�>���r�`�͖�Ѕ�V� Kv5��iΞ�kW��JA�r� $}���Ӷ%�u����M��*�93�q�Th*K��>�E�:7u�y��	��G��6��bm�����Uc��!~dv��7�}kw,zuCs��- x&&xhl�~�Og1D݌42��Id�G���P��<�	�#G��S�[�fOG�H��f�x�~AH̷�V�XƩO'E������bA�褍�ʝ4�+���4��o,��M	����v�0�����fH��ଌ�?j�v�/J;_u.P��]S�ݷ[Un����C(��k3�+]�H�@ 4]��zʦ�D��ԇ������	]���}{�VdW}qM����	d���������Re�����{*+uM���R�JwU(�9\��`Q��HZ�[G.��K��v,%=,۬ڽX(�#d���w
���尺3>Zh��y��s�����뎔V`ևo��IQ��N�������T#<S�xF��X�%Ɨ�̣z�[���R��8�#�Y8�l�ի���?EN fvF�}��T� ���r?��7���AT켥] \��8��&��_\M_��w2�ȝ�!i��wr�`"׎�T����GD��q�#!�%��0h �S��w�vA��B�OK;�d8��n�u��*�b#ewI�a�r����+o�(�^��ͬ�"��s��
h=
�	�<5	�BĻ�yD$�֩�?�S�$	C�D?�x�$�GV�%�!����'\�a���J~4�5�zs`r�/ەQ��2���`n����À����{5��nM��'�!�`9�!�4s�w���>��jV��\��������K0#p{v"�qD3�;z�) �.t���t���ǸM��L+Jd����\@�b�G��{	Bmk����&���C��1_�����鯡%�N
��p��;�� �2�%�YܰĤh�LZM_4�g�}��
|j���3: �)7D_��;~1R9jO�' �#l\�\Dj9�/+&J�/��׽i��Y�V;?�����cO�mC8{>��6Rx�$s�����8�|=Ug�uN��6��W��:��/��@Fvp2帲Wg��Ƞ��4�\s�f����I|q�+: �7����W:)�\>��j��ܵ;�IG?�
o.��p�ƞ��\$���?��6Qظ�Jn4��D��4�5Y�$��;�'?n`��bd�h�)�Z\�Ipѕ;�#�k�A������;�pox�M��E��!�0I,"�u�2�f����L�}b+a|����0\:Y- f�2i�FW9�h�T��ޫ��d18͵�B@B�x���<)˴�ybfa׶s����������ܩ��$���t�1�IM1xd:�3���6s� 7�0�b�Z��s�`熈�E/���`͡ANt�ց����X����V=���5�ַ�cuwjޤa���,�$�h�d��Vz��N�������HUv� 5�@1�����tn�`N��+YWQ��^Mź��j�^q�5h��)�
���V~s��D���l�	�8l�����`i�F%�x��h����N�ϽBzA�[�F����t;>��gW�E-�N*I�|�0<w�V�ڋ�Oݐ�iP�Q��^�D�b[gLyo�n��!�$���
?���U_)|�6��R�4����e�d�,��;M>KIoA�L��R�Q6V��C�5L�؊��x�b�,aqb������f��� ΜcWv�K��yDL�[����z)[��E!=ĉ��&Y>K%� �(��-�	t?�
+T��@<E ��������+X��)�`W���g��'RG[��ߞ���	'�lx���5��l�B)��lѿ�;��#$�,���a�3:jq�=!1K�6*f��"px�|Zřxa���{#�/(T�o���x��l������Nk�2���]���Y-(�	�r�L<7	���TS Oh/��ab���7�Q��`I��F܇(v��=�/����]�;�N��L�۰[��&�p�D� �p�@�|����o�r�&��e���h�ҽ��D!�l�G=�� �wG+����4�� ܰƺ0�~-gIHX�\�&��Pc�!VD�m��<q�t�Ta%�hcPm�]�3�k{Ғ�/)Quh2�6s���z�#�"���_���䫱�%�$ڷmby��D��0Kj�d�qlV�C"I:��U(R3��RJ@�M�H��hg|����%���/�4W	�����-0��'�)����)�:��`DǕ���$�)�s�x@@ѕ�/W�����^Da����D�Qc�p�����x\}��H��1�
���+
�����$D�D��Hb�j.O�C
��ɨ����/�`�i���T�)��d���3��Jn�� }����4����� �L+*(W;��| #�&u<~�d\�	��%4_�� $�$�в��J����M�������O���1y�X��k`�P����|Mաɇ�Q諒��gG�6��Yz��;���oՠ�`buׁj�B��7�
|n�~�F-K*�\��k@pT�/DK�W��*�����X4(�+�v(�K��O���z��b�u���<6�3}��n��a�����?���մտ���-4��#K���i�N��6O���M=�F=t/�;�!�[O�X�>�\�[ؓ(�׵�]�fF� �{0�E+��Eu�Z9���e��.p=9Kc������9TN�2�#����~F ,��U�w��kN!���5�J�-q'B8�9En]>frr)a��=��}GQ���.�S8o��=:-^��ô� �hڟ����й��DP��&�9�E�nBkMЀd�+nE��'85��x����T@��G�U��vu�K���T.�d�����C������ѽ.�v����T;����`>�� �ğ������0l�ş\c9���B��S7��ik���W�KZ�e�Fi�/9�><�c�\h{���،�T�Y�"}�_���@�;�����:���[�����m���iM���^�G��E �z7�T*^�"��M6_�A�O�*��=�.�钱�v]`���Iq����м��+�^<8�i6���������윧�C,�e�r�R��~�|d^:�s�����/�-���^55-GަV�]봒<7+	�K=�pe����R��/�̨4ˋ�z�{x����	�.�X0n5��Ͽ 18"Խ���A����v��0�~�Dȧ�B�^8���Dt�q���.��>mȕ����>�a�i�j��c�
�����Y�X�)w�)W�T�<Ͱ�k���gon�لYf�qf�׺ѻ�,-�z��Z�Ǿ��̩$�~F"
��$�z.�/��S�)�6Yi���L�kN���?���2�R��+V}Un^SYO����p `���Ћ�󒌭�n?�:{���u���1F(��˾��/k����3�]�R���Lzz;2�:��T�l@�ʩ�\��HyQ��@v��կ�K�&�z���k�x>о�>�y��v�פ���n쁾P6��K�O�_V�����o�,ZM!�CQI�s���������"�bS_S�!Aq���ǎ��^�Y[�W��PɃj�On���3�D^M���7ǗE˸Q�'��F/<5�%��\�pz��r�u�����i��m���F��.ᲇ�wX��@1�3��p��{�vs>D�/�!U�a��5+6o��`G���� /��H���L�TN��>�����bV��R@���xGԝ�X���)���A ���p��j3����Ku4�/��>�M���d�n`[2��E�<îw�����g줺=ٜA�[N�)��`���Nz�p�O���<�j�:�f�I�g!�=:�췮DX|��R!t��G�<�߉�շ>@���2�R�e��o��B�+�6�qG&,�����H(_M9��E���Z�_kfֿ�uo��@���hsE2/�\V�7�*Tg�;�"/��D�U��--+�g���9����s�:��im�[܍@!B=�K>"�j<-����r���N8P����}�H}�ݹ_P�X9�����_hӫy��_j<����FҲ��'��U	�)>�D�L��(��I���u F�0����*���X"_����-aZ]������/�/�[�Q\@��ǎ�(�l��z>`��ԁ+��닰��B��g	�1:�����uŦ<J {�˪ �*��Z�]��CL��g��X���b�9��ϲ	�&����QGEn�/[�r���B��q+|����
��rxg�M������K�3�=�lT X!<
�T[�D�q����^�jU�Y&��=�O?e���;����+��cnp8Q��߽0�D�->��ڊ+_��q�/�0��I�5',6@&����ĭ���4�;�Jb���~)�Ă4^Hj������d�H��QG Q���9I�￢H��@��ψ�N�b���UQS��H�
36���pbݩ<lsIf�h�G�r!x�%�t�������}6�	�M]��ɹC��M���c�`��8-�x"�T�܅ut�x�L�=߃��5,/�#����}묢��C��;�+�,��;O��&z��)q���V!i�nd'�M
�i� ���E�J1�)=< w���Ѷ�&����	�c��^�\���T�ǫv"�Q�;���4�}����25Kݺ#V ��K�nj-U3�=�.}�c�=���}���plz��9;7~$*r�&D��΄�x��Ѡ�L��_.
��%��̓\��f����2�n��HB�)a������Z�-#�G\�s*:�<�Ә�Ο�9��"J�8b��e��|��{�i?UXBp��'�@���ST��[c��ڇIFo�FVp;��u]J�5����-���(+����$
�����QG��w�hM���o��)�N�<D8m����ڤ���]_A�\4���x��W��@ &4u�JӀ'dV��ۚ��2�mY3 �`#7��*t:3�ψ�|���'v��͎��գ��e4�!��bO��F�<�S��X�w7f{�;�>�JG5�_��n��7Ǽ�q�x~�X~�C�\je)�_�:"���%��1���t��:�����,f8�g����Y��lZ�Mgcr�\ʆg�mզ�ܵ��X��%�W_�܊$z�J���L-E�?M�(mZ�(393��;n���#7�P��ah������w���c���܎�ٝ�U�'_kZ�ٍ_-���q�Gr�5Ǩ̸Nx��]d��} �U�+���1��>+�M�\�z�)�/*a���ޞ5Ω���.?`��(G�dG+�
�9��~���a~���-lW����͌����w7�D�3���C�{��0��&���`F*Kz_��V�l�S������m�=���a�����S�q�x�Ʃ<f$�%?SD(}��+7��t��)��2h�w���G9+�.)_}&$Y�ˈ���E�s��󰗌^�s��!��z�x^Ͱ`��'�r���K��� �Y?�;�5p�3c�!H�A?�(a���n��V��&�l�k/��aMkʷ�����D!��^�*�z�c�,ڲU�0P��$�
΢!�'>��u��X�k�U}Y��W�7�A��9��Ԟ.��J�vɂ��)k���,�{8��V�ޝ@�Vg�Q����@����b����?��{X�CBI���w�[뱎� �B�B�{YT����xؙ�8��7��-j�;�U�ʳ^������]�r�(�>����%�a�g����7�s���k%�,�V[�C�)�	��u)��Go��i��dbj}n�9��n�$�!$�Н�'Rvp����FL����ܱ	�v�y�s8۩9j�w��*^U�x�����7�_Zѵ���Gk Ĵ�ȜP����̾���b7Z�;�s�)�Rí!���h����+��|lP��$���'�2��뭖�*�&:���h/�l7������<Tl�o�>3W��[���r9,��9�'1�s65�_�ޢ.EہI��b�S �}�B�.����dV��KhVj��N�n�\�X*[�IgLr����n�{���.د6����W�_:2Y�U+�&2	[o����}<	�<��GOJ����<��+No��"�d�唓�Z�"�(���Ne"y���pɰ�~��严4І�X��@��[hwZ�?pۆ�m̷����o\�W*�W0a��0�)�����KCl2� ̏R�U��s�����yl�m۸F�~����"We1s�e*��>O[��6�S<|��m��㱧\�\p��/�V����YՏJ�gm�XV�"ѳ�^��P��F9H ��W�j�_�ӱ��0l������g����%�t��礓%�f2#��Y�a���_zD�*TdJ-t����ﺑ���<��
��!|����j�Ԛw�0U~35,��É������w�|��F��k��ې�����l�C�I����[���R8<
�a��r����
.��Эvf��B���`_��}��͟����ވ�YX9QA��0�U= 	�Pl��4�3���6��D��04�u�-���׌�b��8���j1��@[=�ʃ4R\!X���]9��iم�H����YʌYf#@��%F�s`\U�6��m�C\嵫vmc�ˠ-}TX�����&�(��*��;*, �5��.��(1��$�t0T��&(ELa9�����;� !*���"4���0���I�{�V�8E.P� ��=x+푙��^�(q�0q&m����C]�����B�1���N}��A�Y".[uֆ�dy"x��+�u�iІ6���捶��B�CLzk�v��`M3w����ůjI��F��_�
/&:�NsK��Z�SX1��4Z�~c�}!۽�9�P��1�`B�(S,��e����h'��������
��|�sQ����OdPc�,�[\�fx�V@٪��-Z�a�o���a�������
�-I`cO[�O�2P��o���V���х�1��њh����(�m;��al?��>�����i�B�Lc�� �VKWi��=��%̘>�~��fF}���g��*:<b�Ί��v���C�<�G׮����U�u=<���n$���[b/���U|p�
�3�Ւ
TY]`�1�.A��Y����Ҹ�'����ҩ�����
|6Wt�v}�R�M+�y`0,b�~�^���T$�FUH3d�nS�_�Y��^2o�ՃZS{��>���KO����7?qQ|#i ��#��/ �wH�D�C�ghz�=E?%A��?���N��T'���Z�}R��c�������R�S�#�+�mN��m"N�%W��L�WP@����8-�	��p�����X�
��}?jȽQ8lֱ��f)���?q��n��x�=X����P����NK��P.ׯLZ-��I��j	X�W��ވI��_��}iJ�_{Y*��\��W�L�D0�<o}\a�^�_��
~4�O�̙ۘ��'>��U�����a��捳W�?�J!�X�5�L�;[³ǾKu������x����k]�%�1��5�MQJs�*�8��Ϲ��A\���*B��Ɓ�����m�(�&�����l6�Y�)�iBA�g�F]���)�eI%܊��8���U�H�������Yn��-*Y�XN��c%5����*����;�1S9Ur���PPg�I��@��%�!����N�J�CC��t|R����ڙ����]ߌ���[�G�Ӱq3��׺0PP01���׃�DEZ�c	nR����%&C��2#/�tM�������Z���/BʜR'�a��^2��y�{�����)K�|�*�T�'�0�>��l�������<6�w!<z����{��j�sA�L6��^�ă��_Pd���W�GzW��\]�,�#V����6L�J�}��i"7#ü}���d��#�ٶ�_E'�+ނh�e=���UM���j�茇Wp`8����rW�jǆ�ץ`R�:Q��ĩA�|��%Wvd<�1�C ��,����r�1��L�H*}�<7�9+��(�R�Н솀�Cm7������o�ڌ��?�l��_E�2u�9�ۢ����Ⱜ���d_e���8�3d�/��I;jP`!��e�ThN c�5��i���N��%|��t��R�������lg���C���e�N�@�ҫ�dH��PtL�l��B�)���z ���}e~���̠!?��a���T3���=�����r��O��n�W�î�#5C@�w̚��U�"��;#�d��'$8?]�Q��8P����e�|�q������fwA�2�m���	g05�^@|0�M�)�.���K���*�Gz���ZѪLz���B��N�[Q�h7�%�1@������$�N��vd�zm͟��/
\Yjd1��E�_�ݰW�Y��G�H� ��1��P�r}�1��hA�2�!��鑚��Qs`��m���8��B��CLM��#f����v�v+��rM���p�u��:�8�K�O�Im��m��t��j��oO~~P])˝J�ڨ�/1Va��; C���w�#v&DL�|5k9� ��^^
�>�����SԷ����l��3SU�0����cI8)���ߔ�.ʬ�LG�s��G�馒�u���G��8l
zHFE!� �bdS��O�]o�B��/~�}b*	�����y�Em�c^�:�-�}�<�/h6i�ˢPY�Rڵ_K_����8�`��|����P�bN���D�L��ib��dQ�0����'�q�!�ZQy�t_�th{������6���a�}�I�����I.a<'򡾌#o�u��h$I���5�639�_h�s���X���r4�y�$P�g�080�l�6r*ݰ�#���U}�:�{BԎӺ�����n2�� �_�qǭˋeDV�p1j���dm��_�/�Z������2;��,&aY��\����n��s�t��]�����|c*Q�M?���@�f�8��9b�x!V�>p_ZU��<�h��ZWm_��%z��������ٸH��;���u�;��%��@	�>���5{���*�K��E�Kvw��'��o������)O|����m�:ڼ~����!���ǥ�Y[аU*O{`����**��L�6^������_J��,�ꬉGP���Ǎ�_KH�%�cX�M��`��Y����Fhg�wq��X�ƍB�橄�.g|���b0^�,S$���@��t��G�i�b�Wc��i+ߩj��.Zf/��4�c٨��w�Y�?�22
mr=X�<JC�(���v��EҢ�!|����Y+O����?:_|k��記��b�3���2U�z�	/J����.��7���s���^؇����kUϱjGKE�M�&�}ӎ��_��!}[\�� i:��6�a��S����06�I�g1I�^�@��ɑ�b�6m�ĸ�W?����e!�����^�^�"�4�a�u}���������iS��@�]o�Ӂ?�dP�UMU�-x�&�lȽǟ�2�;�������mMd��%�ߥ�z�[6P���x�s�	�Gj�va���ٮ��fE¨��D|���{�d�E���@����|l��[�L�md�q��e7L"E������N����kQWf�E�4�"��˂PEϪ���C$�؄�%T��X���֑~�0��e�/�g��vy �rR[vp7Iv��h��-�fp'�Gx-�Y�d���%n��������E�����V�d���n�z���wߘC�����5� 8o0%T+�B`PAh�K��2�C!���A���P�5�������A�RrP͐+)�̝n�@C'"^�Lϋ V�QF��F!�:�|%aŭr\��Aצb������L$;;����(����A	R����=Iꔢ��j�{�A"�d&�*h`��rA�2�{;Đ�k.0Ce�˸m>LeA6gd��X<8��*��aK�[@9D� gR�A;,S
4���n<�z���<�V�ŵ��E8):����$U0��U~�P���b-�K�C�m�$f��,^#�y����M��yk�d���h�q(@�-���������'�Ep��$�Nn�Okh����ɘ�����?Em��7�H�^�� )m����n@� �H7�D]	SU��m�VN�IU�n����67V��%k~.�Ʉh�������࿑����Wn�jS�ĉ0��Q:5�׵�����?��z� R
����ݔt,��DwG��w��i[������'�J�|%\�$+*��ft�5X�6:��07��;&�i�>f�ƣ�+�M�.u��12e����;�~jAD����'�*Z�d�J�$F�7�Ev�@�@K��J��+}��W�Pͣ��a	�3YP�K ����5'C4ʘ
2��[@�}���*�=�'��ŏ6p���Vw���Seu6r��3�%��xt�rh��G߹��j�v��,��6ȧҡ-xD�V�w��z��|K��F���r�4I��X4�۩��x�
��9�h] ,���hz�`�U��p?&��6wQ�#�~ɦ۫����~~�e�t�R�f� ��i����A� M9h3�Y$Qz���R��g�:�9�'�V�q�3���`�I�U�h�����$ܿU�1����3�.~�}�P������Aɰ#�p�6ࡸz���n��XءN��!�K�	{@f���s�!�bS?x�ib��� ����G/&�э=	1�b��dy�d-��kn�<�:��BHP�ڑR@��� �H]��/_��ǎ��<�C"�EB!a�I�/�h�_w�q���P�y��P�CK=�:����͇r[Sw��ńtG�Q���I[�!�$�b�/�	f�/*y�˾��/��2l�G��@d�l��3�pi]7٫pk�$�h�w�T�;�m��Ď�#E��ւ�`>��ܓ�o�d��'-�W�:7���!�K�s�o���K�a������=�����q����1k&��V
�J�x��&C���F���� ^�M�W��曽�D�W�>�&l_�����eXiIowI�]-Ũ�����d�T~��>��t7�������������]�3�km����/Á���9c�tN�+*�*v�'���\�{&�_ Gq��2��끫�y�<[2I
�s�r��S�m���g��E��7�%��_���|��ϡ�W�^��6��.��b$�T���1T�R!
�<�������[���p�)��]�-�H��;W�����
/C�����"�ƈIo�=��Ҫ D8H�5������k�3^a����S�X��J�y�V�TJ����J}��9B}ﺗ�O�dߡ@?~�u�����h�$p�Y7� �s9���+�!%P)U��M���1"��u�rC��~:�3�44{$m5ČC�aH����hKmd��(�2�N�RΥj�;i��8�}/ө���=�&�a�K͜E��?�"�dh���F���p�� ����H1��ܪrcL�5S˄_u������G6�\g)�	�pP\��K�j�݊9�L��'G�N��j���~>�b���q�3�h���-r����FH� yy2��?B�?���"�߮����}#�j��0֫u�*�q�v3up�Y��=B#F��5�V�A	��~����u��<�Z�{�]��=��}�`�ڂ�|���ݠ�o?M�*������OںA1��|�������w�	�f��"���`3��7!1a��=�f��@��L<艆�2?n�����B���/m�x�e�B����2O��M�G���7Z]#�|-�л� ���B>fL���h�x�F!Ê�Ŭ���t�AI)ڕo �F�w$������T��B���/Y��5��ܪSz�X�Ah�5�2�tcWȳ?:��K��..`�8�L�dJ"Ų���p���>����]۸��K�r�l�����1[R�fv���WŦ�$I]��h���#e}���D�p��z��� [��-���h����d3��=W���)Fv�Ö��U,]����XH��������&A;��H����>1�!� .�#�'%��a��3����	h����K��ĩL������C������vT�1���U�i�_�/�Sm����z������	ۀ"!�ޏcp��ܽ� �^$�4L2K�X��6es�TIJ�IX���W3�`�o�o�cM秨fԚ@HD��2���0\���͵r�_�5���3��/HH��z�g�J4'��O_V�{PjQ���0�	�%i�Sz���_��k�@/����]%��VWS��=6��cu��� �.�Լ>{��&�(�ΉT*������
n�h��G�0kj�iS���kE�J���������df�ǧM�������3Z���iKH�[�{�5w;���ӽ�ey��ԟDkC�������b�L����N� qΚ0��NW�3g�H�`�@�T���[��}+��&�L ��� Լ6�ဩA�Eҏ{"F�z���`V���e'�&�lTJ�~�X/\�r^2��h��ɟǑ�C*M|�0/)����v�,'.���	"������bd{��H��m��@Ց}u�r��fY b����?u{�DHv܋�֍ɂ���˱����5h�͍L8�'3�9�Ę.6�'9%4�;+�;v#�qxX���پ���> ��W�
�=K��ɉ��d&����<O�+m� _�=�aZ��:^q��Wj��n����������cDw�{��N�#��͎�c�~��/ �h���;Bv���(�(�p%�PQ�I���������|���;�c����[�g_����`"/��n��ybj�nس���zXu�۽&.�.�P�ZuG�y�)�2!��E�ֽN�['���O����&ّ7�����<l���F,N"���Z@͘4�y�R~5)M��k�3yhq�pR�D�����If9���*ߥ�����#���³��c�y���Hp}�+���6o��zݤp`���xnJaO  %�<�>i3�F��Q�A�$#��%��k-lp�k�9[�Zl��e��[GP��i��P۝?+�(x!����2p�}���	�z�8z%Q�h���|О�YZ��A��By��[�yxcƶ�}��N݈vu�[�Le��Ѵ��#�����נ��1�yĠO�Nm߿9�H.g����'����M��I�M��}�œ˻��7��G�
fsv�/��p�W�6���N�i+�0��Q`3''+�QBRY"}���#AX�Ր�CC`U�s��o7�VŁ�_�Z�\�A�5��%y
[�����!���M�kz�fT�К]~5��Y:��+�D���!m�{��b���?5f#��Wp���[��ŋ`���.B�[!"�ާ%?r��;�$�۳�=.����`�>�K���&��R{2����db{�mkA���@�-���&N�{�rAMۧ�.+l�u���5��] A� �$����{F]����\�r�'B{Z�5�pT�a����Ǚ����h�KLh�@�Nbi���9�C�h�8�?��B#g@����d��[n��������F�MH��i3��@R��G��v�˯�z�,x��E��FZi�Q:2&#�,�L�)�wT�ggEM��z�dF^~��_��m��b��'����7m@��j$6��G�l�z@��怣�:T&���h��D#T�Ҙ􆗐v����<��?A��bq\��-��PU�ڪS�:\�ضI��4���Ti���ʊ�`�p2dq4d�����u�i���F��� ��^:u�l�v�9��yR`�,��I��z�,)����kBj���@�6��I`%k�����|�U����խwD�ٙ� :���gn�<����(�mWoA,�.�H��P\���M�[�����0}�3��Х�j�0����n�̐Iݭ�'ê���z�d�r��&	#�W���X��!1P�q��κ�`gR7��v�0�!��*�@�	�:#Ɖws*���-��ǜBZ3� ���E�2S5�h�ˣ�H���#_����,���-�+@�QӐx�$����c��
O����}C0ʤHQ?(�61�ӍC��T�?a��el�)BP�����9�>��ڴ������t��]�j��YD��v��*���+C�����d���f������K㙇��d�珟�(>)�!YҪN���ePs�����/��
�L�𠐇#J��$k����Ƴ֭�1A�=����HU���&.�}s}sֽ�d����,$G� �	|�HxY^���s/�,��'��|��D�B���B|��/��"���2��և��A��i�)�F�+��}d*�	�I���&ܭd��gHTb�Am���l�[I�%�\u�pF
f�V:s�6���-�ౠ��{'W���w��:��3�4@�n���	(�Μ���z�7u���Dc�{�8\8G��Q[��!+,�n�Q-4�#{3�HUM���:=���M��X���Ω��K���ý�MB��:�j�K�)��3)�/������<�����xQ� dwk���x�:w�����kc��"�y�T���4s��*9p�Gy(�zC�1��w.}��Ͱ������d���#�^6f*'�C\.rn�m0��0[Y���s3ɇ�q��OSm�1�ה2�>}�BKre���)�Y%ʚ<v2/E�����3?��d��p�P��������-h�q_�JQ�Q+�b��Oj� S ��m������=F�3%}y}����g{{$���JEE��U7�_��X�JyL�a\��zm1-5��]�;-e[s�g6{?qԵ�E���0
�Y�踃F��x�
:&�����,λs�a鷭��B�M��2ԊCa�l�v�������ܩ]��"r��l]|"j�Kp��܏��n����h����
��+�v�F(P�+���:��!~�W�z�j�
�ъ��E����U��}�\D�1C�_��nt�h5axN���C���R��|�!�!�ֆnm��Q�X�m4n$$>krI����J��4��z�fm�/��'fD&y�� ���[5��p+{�3x����a�D9�=��]T»QD>�45��G6J��BHI�Ȕ�"mʛp���<^ ������j�����QO�0��U5v�}4���ї�N锋�V[(�e��tx� ��A*-�i�l���l���Kq�D�j�?�Z�L�v[���|���4��$������ ���S�Q�ϴ�J\԰l|c����bMl:��.�3x�����Q� FK��y2� .�Oi7��U�}B�$����Հ0��j����j  �/z�iu��e/�~����Ï�&H*�:�M *#{@�#&F�����/��Z�O;� 5ZN���o�k��O�a�E����zbw�ܽ!%O}[ 4
�P�9c�����UҠ��"�i���a�[��0D�c�9O��ę�dZT R]ץA�&�\�ɑ��As|�s�30���-4��yz%�8XU��q�A��G$�O��
�J�:�[�c�e����>�
U��g����Q����%38�F>��ݽz�i`��#	��.�2)�Z��?���a�EzO����^<p���H [zw\�W��%{y��f�� ͧ%���E��6�ǔ�\�M��1O�����)�Z��U�� $��Z�Q Nn8�Ƕ=�k���}E�,.��9T5o�0�����b"�1�9!�nT�YOT툒U�N��� ��f�a9M�F���t�S'���BnX�;uI�;)x<��ש~W��$JMF�oM"�����ޫ�8+�9a/*��m�n����͊ -��2ro[��"��qE��aV�_*�  na%�|R�����l��F~��D�f�AN�dl��(�����2A}�7�Soׄ�X9����K.�C�
g����~<M+�Ƭ\�T��v�!�6&��ӑ����|�P�]�)��I[�-^@��������x��H3Hؘ���R��7��� y��kR�L��%����Jc^�nQM���ܬV�kC+L�-�Z�5�9gfB��oZ�ZJk���#E��3�o�ߠ� &���y����)�&���
�w�o���F���������1y�xi歱�+����Ɓ�h~�oqC��v,Qm\��:�,�^�,�����T[�T��fϮ�NHL|�SH�6�!��3[Q븩�'GO���^���me:�$2E��I9�����?g,���
x+�ZA�O��+l���i��E�
QueC%fO�������T��4K�8P��m�<]�����L9����`��q�S���)���:)��u�xg�Dٴ���0�/�z�'���L5��yz $N4��W�A�7�X�{Ե�#�ĸV�MJ{>A-�&�O��C�H�	6p[� ����w�~�R:&�[�������U� �ȴ�Đ�en� �`�[�WK�#u���Ѥp�E�ܔ�	�K�s[;/�MӀ�	+(&���\�Yz�r�Wr*eMLЂ5%��zQ�3jU��ke��Gw�$�١,��mƦ�Sf��jt)p?<����V.�}HI�hpQz�2��y$h�W��%w�,,�^܁5�)�I��+���
���kpN���O�guT4�|�Dt�3y��I:����cRƢQ]��z׿�ҜA|G��`��U/���f���w����F�nJ]��D	���Ejeg��Ҩ%�e0(>��M��Tf�N���rB��pr�5@Y_*��Y[`��rv�R:SC ,�o!��0��Ryķ������V_Y	k��x����fH9?�
��ms�7�K���O��H������r�Z�Qy�ir9s�,ϔ��]���Y����E��Է :J��q��7%sV�S�҇�Q���+�j�l��Z�c7?������[-��1��� �W���Wun9�z~���~urlMY�&�O�c���L��E�4*ۯ�%��=~t*V"h����G����h�]@ �ˍX�'�9N�4�a��h"������6=[o:J��Z���82W��M���vl*
u<��e�b(IN[�̼p�O�O�qJ��ІO�dw��ʸ�i"b�+-�ۋ(�fTLJ2{�ɑ7�G���i�?�%Hj�o����]ڶ�U��cw���C }��=z
�\ *�V�w�L��Iˑ{�z�2T��;(�&��t�au*� OlH�
�-�!��7dZ:������ʕ=��cբ)d�G�������2���r���T�����Eۥ����	RC�Nk��#�?/�/���d�u�֑�\��֭ϲsNe� �<�N�ޡ� � Ra� v����g�
GvP�� TV�ڮ�e�F��{!��iT�@���9����f��~͔��T�TA���<�V.�v���=�5��JcdP�Ul(G� ���
�Г��\`��
H����OAS�)����HC�\��J�v#YWc�P��Ґ�c��R�(��gc �6g1����-���L'wב��F6��xxamh=.����Rډ�	�!��ǽ��BF��6Iq����7�ѧ��R(����~o$�W�O>�p��:C�k=Ao��t�d�BB��7��m��I8�#�`���ܟa�c2��P��ᳪ���F�t�h��iϑh�&���v~Xc��SHd�%���A���7�!�o[*N~*6Y'�DD�)��)7a"_���.��:7�w�Qe��`��{hk'�"PK7�zp��쑂����gr�PE��.+�g�߬��r�����D��K���i1#� xH:�2ct����ǋ�"Fp�&u�X9��1����d�,�/����jUI}�Ƅ�z&� �]ݡ-�͋���� ��:�Q�b��F�2f���*������ Jak���.ON);����VR����-T�	 ZS���ԍ���(�x�b�AR��ݲ�,\J	��2]����"\����JN(�R�b&�j!�{�Rg 4A��8l�	@X�����d�u���"9��UIC����Cf�̴�h�j��.��V�׿��^���ſ����i���rzP~��}���b�gsV��C��\D��v���ԅ�U�.��H���R����6,׸@!���{X�Tf��#�_y��a1*����P�1�"��R`�ha�P2p�\Swċ��]9�]K��(�Z�+B��f.
6B��6*�_w�1�2$��N^ZW�ǖ>�մ��!S��LR硶� �G����������RE�Z+�U�G<�MC�q���z�޹��x��f�3�ۧl�I2~���3�k�G9ȿN���ð���5�;?�rJ�މX� -�.��I�Ϭ�O-��0� �k��H0�x����ֵ�����tS�I� *:��Хgg�P��Jz�����/��IZR�`z�0y���1-(R�}!�F���C��R�	J��s?����������[���G�������zH�u�ܐ�V�Dw���lT+L��
�^^x���:��|$�`_�x��@�i�ǚ�ԍ1�{w �C,�Y.�ިZ]�V����(u����r]�	>��S���L���K��M���	6Waơ��>��D���3	�e04���[^�mP����Ο���w8DjE�����<�L |�DS���}���7y/�+]�ʋ��e����"�'�o���Y�mqN�������cX�~��&�Y����?)����:��&��r�l��<�ڽ�"H
\���<;��Ag�	��]���E��S4�4wH��.=[�#O��$�T�zp��ep�{����N��L�M��Wr`�u��b�J��w�<�}�]z#�W�+.�ś�Us�_}&�p��؉p����X]VÍV��%���ot��d��t���5�܂;�9�����m"��R�rgӰ���uBÕ��óJ������:&���D�'��#R�l˽k-
�CkԈ��s�6�y�R�K�B��:>���j�t���WjۚE)'�����I.%g�9'����棜br����:H�-�����a���%��0զZ�T�ǥ�
b;�܇��?�6��մ��H~����\b���Բ�5�b��z�IbCnɚ�'�yN����P���"�R*E�Kv��fIfɸ%�����M,dJ�W�Q�� �[�L1Z� v��Jh-�̳�S�Y�jK����b�4���[!���E`z-��}u�X����ǹ�w�R�*��\rV��x��l�7��t�#���:�l@SՙdXzV�ׅr�q��J<я���^G�7+��F"����`�N�R�=^��o>��6��z^1�:<�׽#�v���-r��q��(0l8c��.��Q%_��H�Ѐdf�����8d;�?�0�>׆��Wl\�x{V��K���#���@�	�NH��u�T�>?��1�Z�Gdh}����U�aU�Zc7O��vGa2�W����ޕ��w����K�Hm��Z���9�4�5m�������Ȥ�F
�\߳O�8+A��&5Vd�q��,}��E�R�>�KR,w[�T���1_-��5,�<g
������� �S��u7}�GSaU/
���`����5������k�\p�����0�����g����m�Q����*�hĞ� A�蔇�2ǲe[�x�A�U��tv(�W+s삡��=���qy�iT1��V���2M���J/�GN�[����e��q���K��!jIe��\�K|��*�`w�,/��J�0�xA[�� �q�{E�6I�E�tAľ�\A���!r�{\8�&=�Ȉv03���x����Ӎ��|�����d��We�Q³���b�6���2+';���=��2�-���GJܼ�xs�C��*��ғ�i�$D�/�p
mSȢo�����-��0+�&�3��h���T������A�A���.+>���p��Q�.��z�<�[Zs�b/=��g�X^����$�v[P�9J=��C�h�+f��ښ����m���ߥ�v��t�*A〲?x��ݚ <2�m$��v�c'�T��y	�0�����-��������i�E�Z̬6�9�/@W��.�-1 �U��bz���QR1^�u!gE�h�%Ϡ��#�ޭ�WXXbV<�5d��켔L��G�Hf�5�;_j�L��F� Opȯ��T'�2��`��"¹�r-�������[U�IH4"z�L�阴�\��lK	���H+>��
�Z�R	�=���vq'i���.���kx��w�zy�
��+�����/�0�E�8�13�]vv��o���[+��b�m�܎�����Q*"�*a&^YW�]9o�]sy�]x��Rh�E�k2Sh7/�t����)۔\�xg��B*�$�K��=��Ηl�����C�Z�U F�V,>���l���F��ٚ6���L����7 �>p6�d́<�s��n�W�P��m�)OJQЉrz��)^�]�>?�E�/W��;F�0�g��s���p;6�)]�	nԣW�^#.��e���7��c��z{��bO������ǔ������Tl�d����SL�+���s=O���bߡ!�e4�0W��Rj�?�6/��2��M�����֭�B�����+��:(����D���?5�W�`�����u���.���<�����w]�`�i�qL�K.[�������n�Jw��錂�)<wL}6��&P��D���j�[ѕ�d�yc8ۡ�LEO�jtL"��8^E�~C�\���S�>z:fLv��u�V���6L]����m���qW5q�/��b�G* ���8o�|��,���u����=�M����?m# 0:��b��Ae�8�O�9��<҃Ab��K�x�:A�ԣ�?	��-�zb��H>mGA�Y5Zcq��7JE
��%!V���G��#��q������!�})���o-wy����*Ӧ���L�vȀy�d6��V��ݹ�Ɓ�^(�P\w9(���%C��Ӄ�NKV:'u�]�ъ�k��U��I�r�B�o�95�?��8�T�P�vB���� ���[�ờ�Q��c���{�W��D�hƑ�����K0�m6�ƃ�Ts�9� ���s�v���n&��9��}/=�n�iL��@.�AQ�.?�)x�S�!�D�vlt���X�����[7��uP�Å�#$^�����b@��� �P<|.�!+j"��CY�i����7��M�WEa���
n�ׯ������2�\�%�ޥ�o�p�dS͜�����DM�'��f$QRg���쉨Z�D�i�,�BG|-/^/1V���o�%4�@�LIi��O\�g���u5�+M�s?��ǸƜ��o X�F{))%�9�3���V^�6ǟp���Rճ>�2��K��F8�Ŷi���Sn�%�w��~ٓ��.!�U��ӳKT�I����}�?���8"��d���Q�/S��}�`#��ˤC��wޱ��^��ո�
ux	wD[x�w�٭3U��ov��G튰*����E�|R�|x�³�A��*`���$VX.�^�S0)*�?@;�_���CH6w�R�fZ8CL���QFE�?�<W�waϑ�.�?�b���W(��J�yѽ��G`>�jfW욧{*�� �B$i	�ʟ�����+�����@�.��Q���!��u6@T��TS�~��R��TE���b����_S�懼#�:#�M�3�I���jv^��	iD�%���Q�����m��j� dN��Hꎏx�/��{��/�:��
�B�K�}�T����Y�.�m�Y(�|ꐅwd�h�E��Rʹ�K%X�34�Y����:t�0�ͭ�5l�g�
����\L��_jD�ȉx�Q[�H9��/��K��[��B_{o��~��J!���>�E�������e�E��U~�a�q�.�o����x�)�b<^��G�I�c�b�l�X^�T�"�0$m-����> ���e�QN��/[,4��7t��e���$Ij��z޺WC��� F��K7	��{���8���K��&�`�D����/�|����������L�)�.��jh�ܤ�B:)'wRrk)=	�o�m�ک��D���t�//s}���|��O�4O�����QpHoVm9�h�Ǯ�/إ\K`g��#=�K��#o�PɻQ־���d;Ȟ��]
R`=���h�N0b�#â�	����_	��=��Y\�ϥ�<i�O/	��β�O�.�^�j&l��G��#���J��78�e�IN:
��M�!p�ށ2s4a�l]�`�s�Lʑ�ڿ�6����e��pľ��1O��5��#�r��H��)��t�i��bv���%�uF����B�l|)g>�I�v�BG�
Q��	y�A���z��u����O%T�g�%�wg�H��}����Η�!`H�`���BQ��q�6?&bx��zC��ZI��he0RB����)&�=&-��&�-g/�'�`���d)x]��Ԥ��Ⱦ]��;�OU��eK#��F�cp2GX�ϳN�9��.f��|b��S�R�M.�.����"(�����Q� |�m�D#��҆���ȓ�d���^���E&d���oR9-o�J�"���mgd����!e4+M�r(�dC���jZR�T*+(����9�-͘(�� p�@%b�:�OJ��
|��^8B���_��3���VD��o�Xf�C����E�	n#�����29�Û�M[�J�i�tze���4��>�|��r:�ywC
��g�%�F�SЌ}c���q�������o.�к��Ҥڝ��d	T�r����}�u��ϒD�MX���F���=�ի+z��F΍Ҫ,\Ѿ���V�+�R�S4�5
f�<��C�b
+��h'N�����B]�";�������U�՞6�֠���iX��05�#=���*��Ȑ	�y_�<��,���8.��Qn2���'���6��S��ߕk�:r�S��s\�M���Α�,�h�=���Jd.Z�R���m�q��2��q��h��,ctfm�1q)���{��s�q<�}��V� ;7�ni��.��4i��72�=�Wt�Ʃ	 ��l�$�u�`�INL�h�m�[��x� ��	�6�w�>g���K'����B�"�������91�W��ӕn󭤒���\��֔W����
�$�$����ed�)���*�"�AZ��OX�XWk�@{�+:J%�!���bH8��2!�R'>�xμ�eI�F�B��3R����"�Hx" X���v׿��J��'R�iv�y��v����X��ī�$�����?z9C$M�[{�%���q��QE�&�De&��� ��Hh���A̞=M�B�͚�X��2����<Sd@���"�R�ߴk�Q`im�OGIu*g1f��bҭ�;#�����Y�Q��- u+_�5K(�۵���5�A��%��"g����!���*[�B��>{�ws��sz*�4��
Czr]���rӑ�6F>��Ta\-�����2p��H��r�eΚ�$=ɉ\#p=,/[���~���¦[�h��C2y7��F� :#ϝ-I�VFP�@�č�~&I�$�QI�TJ��k�Y�	�%�vM'.ia)�<�����TC_�w�!��87=�$��Kv��7��^�'�L�qvCDu�hs�33�!�N���Xg�NK7�+>H�[�[-l�����1�
����/q�:�W���sVV}	�>�C����Fm���3*��A9n4��RcE�(@�r]�W��Q'�?��2dlnBS3�|dT��.�$��S�!�t���f�w�=z��.Q����]��X{>w/�f�?�E��E���P�X�=�u��A��~�Ͱ�)�Z싐R���~Y_�3�
�S3��= ��j�����`�H��\���d�}���,��*m��O�)����{5�X���>�� ��њ��ɝ�K ,�N i"��<�� Y-�@���U�UT]���M��j6(��}@?����F����zJ��M��������N��M/H��hZ��C��/)R>e����k�ԞR����-0]`�\OS����k�_��{�9�_�.��x�q�B�1�k�z~/ɾ:Yi��S�����+���~Mz"y<�����^h�#rBx4���/�=�@L�������B��73�E�w>�	Pͽ?=д(Z��e���z�յ�|�IluQ\L������82��.�`�dV�s�$�xt:��Ъ��l�f���Hi��D,�|���P�K"OǂՉ�s�p��ۂ�J�u��&c����r�\\+ot`��u��a ��2�n�0'�\B�
i��Sc�7ZR�GOo�͹�N�p#�Ѿ�h����c��*�r���r��@Ik���>ڙa݊\�A�W�iM�E=�z��D0��O?����E�][&{>)��)\d�?����[!���I:mk�g"B�S�gp�x��.lBv�I
8+h��|���i�5���2`�E��,*{/��$Ue���N�})���ˍ.��S(�3�b�ǆ�$4���A�xvdh9yLW��7ͪ���3�啲�ӊ��`�+�'oud�4�� s�CO2�NKL<�)�{���W�D'�U$k���6�yn�Z�/%.� �&K0����J���.� �	0xE���M����ʯ�-k�L�U+w���0�>�����/���,������[ �4���s`����X��<�&w����+eb50�לY�L���i&Ζ���ta���������jy��т�z'�L�6�H��}��V�k����
�$ ��y����w$_�E�jBZ7m��ٹ�E��O�'�o6����5�?�A)�����<��"�;�E�Y�Ky�0qj�?�#"�h�#��69U'qt��fv+T�h�a�:�I,���W�I�9��
��L� �����yN�0��*�|BGX7}�������@��z �m~�/���7JfOB�[Á%h��`���L��\��Чp�ٴ��-5��E�Yom��2S?�fW!:\�Y8�,�V��ć�Sp��gq�9�O��}<Eo	�⥮�G�=#t���Oh�����/ �i���S���E|��muu}��lok| =��X>�T�Zݣ]��:�g��j#S�ړ�����"�����G�}�lC�⼰�.��"}�ʀ��(dK�+,�-
�:	ңP�����|ab�1[9t�!#��O��zoER%��?�DBS�lA�!׻��W�b+�Gw"����FUZ�Ƕ�Q|
0��[�
��Гz���#�98b���Uv(��!w��-���p9�h�,ǰ��S�+"��>.����C��f�u�9�>T*�r�l��r�^Q
�5���C^!�Y5Ĕ���X�#�W�߅����}�O�ħd�r}��O0�����R޶r�@�WP��E}ݎ���r���l>;�'r4��5T[f1�lA5o�� ��E�M�sJ3�ۉSK�cJ	z^�Ο�*�*.��_S̡b���0
(�N�l�*t���k��I���{V���� �� f�yaB�Gp/O�B�!�D{��.��2MتS��>w���K\W ��Ӕ��ll�<�U�S��g�.��ZEY�틻`ӳK�^�f����C+_��0э�R�6�!%�?���B]����]):\��/uo�K!����?�������Po���'T�����0�Z�B[M�����[���#���ݚCk<�oО��]�Dtxt���Q��~&��^�N�[ЃWȄ Uy�/~�ae;W�-�`�����HC���|%�Ǔ����n��Ɣh�	Ƒʇ���r����#��#�va�:�X�Y���8B��{M)) ��ߌ��GXɪ��Ʌik�qD. ._,( �X�GIk-��1�f�]�n�6_�%%v�m!a}(���P������#H�����܌�{�뜬�O�1[~���6����9�h���P�Bt�*�9�XB��fH_�o�0@19�Iz�8����R3 +�?b;c��Z&P�w�<*�cj(�n�`�
7�+���$Ӄl��?T��v�1G���K4k��R��Ǉ��Ф^�a����^�G$��R����jW�+�UK.K"��À�߃����xU\�h�Y&�KWuJu�
�P4��S����� 5�#��m�a����yTJ��Kj���C���t�z�֒���a��&��n�ս�͵nѪ��v�2�?,�SVVjuX���\�u��k\�Ш�d���_�N|.3���[:@��t��a��}g�g�����
��,	�<�BV�3f��0�
�G�.6G.�^���ǘ�a|�R��M��7�(6�χH+�M�7��g�hN5�=�ߺs���|R�ƭ�1!��Z����n�o'&��ɫQ�`LӉ����+[����W��U��G�k�%���� ��y�^�̴���{�*�C8�a�r�o�x��"�6�IL�=u"��N�_�l�Qd����PՁ�Q���9yړ3-���5H�LhRi?VK�z�+EI�D�_G��NP^��׻\�{?�r�v�
�e�NH���{<��@�}ߓ���Z��l�x���Fs��N�9�⻫�ɖי���Z����Cǹw��ߘj�˰N�0��+ߎ�\jΜ�19���9��t@�q�W����e��>��a:��K_m���q�o	Y~�\� N�R��S�+�f��ʕ)�.yoQ]3SOQV�*y�[L�=xp=+��2��8�ԡ���c�7�	�[�֐�3�E�,J�5����P�����nx�U��WR"�$��5��}Y-ӭ�l�_}����!F�����TL�'��@�����p&ʌ�en�����'K_�A�Q'����^x�Y��<����d#D�Q��o�qPA&�RI�R�}�&k��p[#�uǨ��ҧ1[k�l%#X�Җ�<7K���`F��m�*@�{��]����Q9�s�K��A(������>��V�׬�����]Y.�NY��R��Uݒ4wX+p�˦ꦉC#�=��U�>�|�ґ��ֺ�����3
U���*)�]0��j��x�6�����]��ǫW�������Z^hd�M�<���8	�x�y#�����&};t�L���3��3\/Q�p����J� �y�����9[����nE�v	EtU���\~��o�8<�a�keW2^�5%S8���mgҡ�a��I����}�^�k%�7%_\,�;i����+P��U�a
"K^ /�PGlU�\~WQW\�T��3BY������<���	Gx�!�g]��i�ů=��nG
L�K8�H�� ��ݢ���gJ ,�e�v��M��� ��e�Q��:��>�tO��gM���H<p�;F�+�`���5��<�1��_c�a1�K��+�c�`-�,�����}�m�<�U�[�� w:�E<ŸŐɔ�`��҇1�q��o#��	����yv�������asK5j�$�,fe��8���A�(�"(sWB?��K�TAȔ<n��f?KDg`S�5o�����S��Vp�gY�$�	��c��G�n�1�xEdz�΅`=���W�\G/u�lI�T�Z�a�6�g����Edzj�E�$��?(�U݃@.���T
�Cl-�߼����J�񧕝ɺ��L�DR)���b�B�I�P���;y���	���r�c��X��Ξփ��jĊ}J'��o+�H'�����D<�j�gj>�:0Q��>v�UW���=�ƈO����M�����Ph-v)<M���`���X�q���g�-7��a��84�l�)+/�_i���q�b���hL/Xa*�n>����)u 	��+ՠy�%~Ф2��)�w�Z�@�gE/�l�I���j��J��Ǳ��">�7/��cS
<���%���J�m%�|����Y�̿`�����ԛ�B����") ��<9�6BA�lnC��I|��#k�g��D��#]�d�ǳ���,���d=�5uf��gn3�ھQ ņ�v���_��*�,Ȉ�_Ώ���R��X�GZ>0V�ApŃ���́�Ӯc�$����Wg��^9F��t���jZ3�aRA��x�9T�@��R�#�c����W�JD�k<o�gj��PH���>4� C�t�����&����[���O�JJ����p6�>�nj��|�A�N�	����d�	����6��@0]Qq����ׅ7�����z1j��<̴�E]:�pL�Wޣ�K �`���Hm�掭Y��eZ,2V�?�BH�{l##���{"��Sv"TѨ7��L�HQ���*i�E�9�-��Y��W���Xi"����ð�d����YC�y�7�q�[���`EO�8(oУ�}g�c����1���n;Bu��Y,=J��뚿%��M�3{�`4E�6��^NG�q�a�� XĪ6̧��4�.D7���B��
��E����v\������ȃ���@���`$�Z�^dۻc$%�,�U���e=�v9���$le�A 3���#��V�OnYZ�WZ����'&(�ḱo��>�����k�Y1F�Na�Z�S������=��T��̼<���]nT�w	"�.5W�o����0e��$>��m?d��@d
O�8	�5�5ז�S�[�qI�R^��}�}��$V�I��L�[������d�#ż1H�6,j�윯@g}����Uh�a�E{2(�Dp��^���X���t��ʡ���N%��1jF�ѓ�:)���}aL�8�>�>�D�u�ɰ!��P�=�|z�î�^E[-@_e��{,�r�F�Q���<� �t�`�J��mV�Rw�:��-5QH���Nw> =f|B���C�Y^U3��55��0˪�^|�%G�(�d���wzs�:�"&e|:���IKv���/�,��4 /��������(5L�ßa�̇2��|3r_��i�Tq��I��sD�8�믻�\�ӓ^ �K���	2�/�#\pN6D����ԣ��֍�4�ح����$;�2����zmW�Z��e/��(��<�5O~� b��$l(�:���)Z�-Ot)2����4,cnH�ڥb'4��QR�:T7����.�/߬=��_��t�ԛU�WY��~f�{3���}���D�H�x�]�2ˑY�o$I����l]��w��x�;�-����h��Ǆ�/��k����ʉ�?��dW�J�X���zݚ0Y��H������t�T@gTb����7�������2�
!a2a��E�������&k�����{����U�9�f��O�^ΥZK�³kS�(x�gꮲ^�)3ڵ͏e
�����[�R4Ѐ ���DY���*P��pVb�V ��Q�'�T��zkF�|/�����X�Ɣ
 �XZ��rr_�kʐ�� xY�T�W� �
�d>��kX�O��Q�|2b�o�Z��E�UFT�'�����{��R��D��V������@�z1R�<�:�<������t�Ғ0T
ːZ�1������2����,b���^��	�a[3��c�~W Dnv;x�w9���5���p%�x,��/7]{ �$��t(K��FCO�#n���	Ip�t�RE��B��Qͧ��b`��Q��N��׀���k�o��}o��)[�Ҿ��#��4�+[�]4�k9�Y"�����Z�g�I�8��l	�H/�m��S��p�t��)	�&1���� <����B�k�;���QMf�L�����.����[�oCf�ڝ�jʂ�����4��4�^#[�����\�ӊ���
5�<̱��z���B�����_u�W��aY}C��a�qh#��٧�u*�=�CR����A�B�9洂����B�]��S	;S��5�6�ei5y]Ě���^�hŽ	"�/�h�� �`�+�wlk��T�Ex�G�2A�\=]��A*�ݹ5�8W�������?�6Ff%c���(�a�h2���a[���S�2�Rк?�] g��{�Q��,n���;�]��"K���~���a���f(��57?�� �Y��gY�*��*�Ų,�Hqz����FV�I�6E��XNS��S{�)P�S��PVHӌ�Pj����;-��e�P���t"Ix%b�n��D�u^U�p����J1�F�u	�ZOk��7H^
�~�V��g�u�m�'7����hLI�⁁!g\-�l�HZv�Q��X���!ѽe�%j��T�bO���W��c�y{�_pN���k.�8
��>��������� 9|[/�d_�%�	5��K���hC��~٭�
��߱�K1���f�	A�S�fF����7�/Fk/z��-�P��+5�~������!�������]��kS��b��	����2��>H�����WU������g'�����F`�ʛBdՔɑۺ�*s��Q�4��ڻ��@�j3�Wh6�H�ܻ�9P	���L�>����;��Pmuԫ��,���M���n���l�O�SE���t@�ȷ��f{R��PBh�	*��4�%L씻o(�/hu9�A%�]�-���td(5A�-A�T�T���a�N�����<*���w�Q������xWU��Ʈ��kTO�#�lK�-��j�
:Գ~#_h�(w���8
�Th��ϳ�5���Is�;���W�/	$�����nF��c�]��lp�K�Fܑ=�u>y%��Al�_D��:���%#K���)��l�d>�A���+>we��G����{�-��&+�k�
{-�p�d�r;�l
N�Ź�O���޻{�q��ԓˀ���Id���V+���n����AQ���[0�0;8t��ckG��뫭%�t�sŚ��c��P4Уi���'�v��W�����iA$r!�Q_JK�gIi�fEu��H4��54>������ؤ�n9��7���r���s���9��@���=�^�Y���U��D4���q0߉��9)r�e^��\�U8��i���@[Ԫ���u�=|��φY{�����Ύ�6@>�$k&H1��]�6KS:���L�?�����8CBm��Ў jE���L�P�T���g-�Z߬Y����pl�����}ߔ���f�}S$ſ��|��A\���b���^�EC2��x�W��c�>G���/�ӣweQHl�_x�;�W�4����Q�gl��Z���E[�C�$�Qe;YcA��3XE�{V�u�v���brj��U�d9����5�)q�'6I"ê݋z��%&C/�{_[�w�����A\];��d�e�dV,��y�=��9����u��K�@��$v�Ń�Y�Q
�._t��#xr΃41>[k���P��ч�Q�ZKz�/;�E�����=_�{f1I�4��Y,�@�^���j�d�y|���r��#lŪ�V�y���_�����$��y���)Q��L�R�|�נ{����L	2�����[͆?��.�AH���)�����CJ������ �x��d��.,�Ny�g�		O���K@1�0A9���������7��(3��*�ԑ�{(�9�����:�K ����L,+���v�&[����'�����E���7�w��YOu�.�c�>b�~�b�Do:h��Br;\�6Yb�o�9�-5 �p+OKO�;W9dj���7�j6_}c�<[Ub�����b{�F��������
� f$��ʯ��zshUS����T)�ŮA�$�L9 -h2�g
o��}�Z^�<�a� ��a����Q2'��y��kz�8�;�4�kT��*��iUկ� �b���_g����
0��%!��Ȫ�hT�c4שּ:-��J��A2|V�����#�,Wf�w�5:��~�nw� �jO
�[�lql�@��L��|���+��`ūx�q�x
ؐF!�6-�<�I v¼@�s"p(A-��|?��c`�Ȧ��xP��M����\�=��/R9:��pk 3�x�E�j���{'
��Y���W0���%=U_��!�ն��}�M86��TfS��'�D��<n<a�3����/|Ϗ���M��=Ƈ>X���@���:�U����H)�7��f.׾l�ڲ>˸~v�"����OCJ]�=����)�+`W�/;��!��$p@a�d3#w&�S4�_���&ӻ0�vL�R?��:z�l��h�v9�t�7�&���R� �"&�����J
�J�̘�y�)w� ���s:��!Ҭ�6�G�����U0F���j��6`�=j��Y���	{3��4�F>�����;���t���LTX)�p��$���"I��f�R��,Δ�܈���W��ٸ7	���u�Ȟ��բY="(����S��n��v��	*��lܛFi��C%���mY/��q��M.�F����ŇdI4�V�4d�����d�ŀ�ɾ�M��{��!�G����R��s��Eo����h��R�nOD}���[d3�T���e��Ne�I��4�!oZ�g��h+/d-�����r�
~5g �'z�o�����Ϋ%�oo ����L+��������`�'�P���w��"�'f8��b�u\� ���	�C��Hiګ*�)���d�	�ȼ��qbR���.H6gw/j��x1����Y3����r���(�h�%�}���ׯ�)���<?U/�'|.����ʻR�A����WG���Sٴڲ{v��w�۱�*����	]����i�汙�!����۾�J�|�����B�cA;��䖈��,u��,(иsIb���RJ����>��T�4�H����> ��7Tn�|e1��i� ���$�dC֮ s�����Xx���`�P%��)V��AɒhBvա!^�����m��"r� `� ��-��rOJ�H�&t�`y�^]�+�c��/�I6o7��?�Z�/3)����ݝ�&���d���y��6�Mrӫ߆}���GR�5mV]�~E��X��u�
��%\Pk�'���KW�'��QP�.��&�/��f��K�u���� \q���?}�&;!��Ǖy�
�,�lw|f�o�Q=�2i�ʤ�F�H��πHOҠE�D/��c�����r9N_�U��]+�C�#%d�����h�&0c��o5�bkrq��j����Q��rP
�o�@o�)Tiy����]�U34�L��������vE2{��U(c8
��gi��>�q�〭�}x+B6�C�B˰�r	;�����8b���lN^���O	�h��&�5�t5��	��������2�+�/��3�]80��,:�koU��j�`_���W��~V����7�!Y��@z�ȰPql�*���W�,㒷�;O�Th��&X�3������p>� �䞪F�(�c��s�)�b���\�� �b#�O�H�T[4C�Y�la�mJu��9���nM�f�6���|�ufXJc��+u�{=T�6|��#�j��}
�hW���URѪ�c$�_��Τ�j��J����?n����zU�%�փ@�Gſ�!�a��/�7"���+[lm��oip�P���]���E��i_�o_&�N�i�����cw��w�t	�iu@�����2?�T	�9�s�z�!�h�x��&�K*GT��.�0-V,P��rܛw���J�DÈ���UT�I
	��Q�_صRN�s����=%����B���Pı� !q��qOe%�Ģ�p[D=��|�ڵ�WRET+�el�j��w��Jqu�}o�{�-^fo��Q��$�5��/�+��c������mԓD�N���K��M7۸�%�'�<�3ndٖ�GԞ�[�^��&Yx�*o������TjF��|���b�)�Y�nv%{T��$�� =Ht���GM� ��q���S���J���25G>�5^�Ѵ��a��>�������o�)	І�t6e+�_��/�k�zG<~�D %�n��2~V⭶�����DxK�˙�����Ԑ�s��Z�*�"��]t�H�e�2�僛.P���I���̬)Y_A鰡�&$�IX#��Q�u���kB�'>iUG�2�22�h�Bl�Q����$���<��B�.��!�
�~7���-bS��e�&�鰁��}(h#��k~�ł�#�թE�����uPdS�*�*!G�w|�l?z�ⱼ1#qYP�&�|���`�Ds��D�[
'���Ϭ��}���ُ'��Q�L
D����.�$ț ;[Q�%��7�낷��%)S,�@G�i��~���c��Q1mnO�KL~�8#@�-W"�R3�kt�����AUЇ�jK֔��>�{U�̀�Mkf�TS���69��a�q�͛X�k�&���?�ݠ��9~"c�,fV����U���6/
�"�;��#SI�8�#{[\��V�;P��=b��Y�IK�=���O�A�'�PE(\#Ը�Ռ64jE��z�}	��mȹ`ɐF�ti�B-�_�8�E@7'�&ӹ��!�'�-/�`po�����0jI�	�6փ��k�'W�n��h���<��0�6P���c�p�-|&�L���
��F���g��y��"��#�y�j���=��q\����V�05�y��쯇�M�vU����J����¦�cCq�\����إ�,����.S�A^�%�M.CF|�V�6XO���� 4;��{ԻW�/r���|
�����,�NP�IϟԀ�.́�_��v��ژx���"r�HQ��rv�}��������$W�p
@mX2�s�:��V�ֆvtr,3�j��1S�[�@ث$��\�h��i���|��m�Knا��6�;�'�i{�0��G2����qrw���ۙ%�
��x �?G� H;�zv�ٍч���8�c0)%$�)��ӂF�^y$U����c���u|��ږP�
�`��$8�gݾ3�޲�|9��?�-;�EC6�%�:G@#h&w?��EB�T N��F���M�RqS�YI=�awte�M¬?�l/�����ҷX~e�Il�)n��?8��>���=�%�hF�����H���?��S����>��-[�S�S��WX�_��3"\�J�=:AD=Ŀ*yfeI��Ld��6f>l��~`~��?�$���l9P^[a�y��M�Gi�!2�ǜ����!�]�rBYoe2iH�_����x��헕�~�j�Up}��ȡۆ�$<����/	���/��u�C������D�>�9��_և8r!Ld�/�
���`l�NU�W5*��^'t���HT�D��/"�/L^6�;b��E5�Y���D!Pb'�6��"}������G�H���{v��֜$.w�tJ����ٮ@Wǩv���H\q�ǿ�����Y�vf�b`-yfY������:*	/���|�����SA�\�3�]-�#�<�0]G�Ţ�<�v��r5�g	��g�Fl�i����su�<��H����_��#`�c�O���^���7����X�OT�P�Z!��_Ӳ/�͛��B�����81˝lq��vC��+�� ƨ��<l��,zWV� |�g���ڲ[���ୀ��Ľ�� �9�˪�G��oq��}��]M�z9C���@n�E7Y-"�.q�_8ǒ�"��3s�%S [�b����u+��J@�r��<��7>�ܷÚ�\5��ɫ-�"��*���ң�{u^�'(�@J<#Q��z^I�]��:�_�m�)��64�i����=�,�����s�V ��Dl��f�~ܘ�lߛWF��]��EOXS�>D��i(�#�^VZ�}p$:��������*��U������py�7�Y��J�4[��|�a޶޻�E��UM���7�������$���wK�x:�!g��M͘�F��f� �PI�1m����G�9o���]�A�E��y]�Ӎ�4�$�f �J��6P��a��q�PD/24�x�%���'��{�`�"W�?���:��;L��	7a�\�i��R9��#�����z���2�	*�qq�ґ:b�V�7r}-c �U�H�:t�H�.���h7�������ܳ�B�[Pz�����1����]`�q�k�l��J�&�Hr�]�t�뎩�(?P��	wU3h,����Z>���)[+��]�!2HO����>a�;L:� ��ni$L7<Z�o��,��nJ��Uq(��b�����(�h@Nsiyy�Z�J�7|z�_������F�A��g0��]��,sǣ�Ġ�^�v50��������zn_b�z��Y�*���ZN>���.F�sL��N ѽy��t�d8u���͖�,ܝ)~M�c��8��iu8�R�d��ye��阀���y��:�.�y�Rw�3W���Խ��s�L��ߙ�Z��g�H�&���r��9��Rf�7����R��r-V�����*���E�Ѳ�b��D����)����*:��|�������^h3D��)���(��[9�5_�{Jw�N�)���cۄ�!2+�@B�N\��T����o��,��KvR�� �.����K���o�M .��;+����KY�b(���_�[��H6�5o����qG0儔rx^I���A��B�r���Ee51 �"6hyA.L~*F�k9St�8UMF�N�@��Xy<y�"��^(6sYFB��*[C]0�Û�A��A�k3=U�û�@�d`���%C�ޢv�+^I��p%�O���<��F��0I�i�rs
!�7Y��^u�Γ,�]+����m�-�r>I4��_M�I�)��g����㟘�Є����w��3)��Z������ �r[�6�t1-��B@��^l\�>�;#Q�J8����@e��d`�)���]��X��`\�o�~���nI
�j�.��S�?��(ڹ��׬�[|�}T��#����#e�G�������5ş�c���G͟,���ؚ��a��mEAT�v�9���m\4Dh22� F�1j�#��pq��V{��˿
�����F2��"�Շ�N�(W�������K�b4�^h�ՆCHb]���;7�.7�K��gxBGB�v*�[�Ѷz��I��E�����z�PAC�_��S��A��*�eeI�֍t>���Ws�k,cdܭ%9�a����[ׁ��_5&��J(���,Ҧ���=�׺ ��~�P��d�t�Zư���Nf�Cg�L?}�[��	=�����gȫ{H����󷿕E�zY"�*Z!�U����Y麃�.z1�?���	����",F���NnbE��yxc�.j��r.��Wa:�P+� ߞ՜�g���Oq�Ԋ�4�[d^�-fS����Dc&G��@��W���f\͹T����,~}��K��C�׆�1ذ
�k7\Iw�4���^�$�6  ��;$ JF�pu@a�ד/���>�uj"k՞ �4-�����������uQA8�:-Fц�Ei��C���})�pz��Z=p�c�1��Qi���,K�z���)Dfa�<�F������$6�^�� U�0�5#��Yg�"�x�7������ߘe��A�����~��zDa�%���/<�4�aA;ٟ�Q�ׯ�k��Z}V�^Go�����������%�;[kp��2N��0r�4Ԥ.zX�c��ތ�E�;]W.���$��7Gp2PFp��;��@��ɏ�ֹ��,#;DU{1Bv��h8�e#cT�%A�u��2;g�ZXdE�xki_ ۑ�+1�=�a���1��E��+��ث{X�qsE�2&�݁]��uTPJ�*�-��7�s�j�r�VMME�|A���t��e=`�`���������?��d�O��/�#CG�R�~��� %�Qm���?>���bMd���$�k��pE�3�����Ϳ���Ƴ�v�c�Z��,��H��� <��z��Ȇ�x�>6�#���ﾱ�Y��W���I4O����V/��w��%q{q".?�V����D��20
Ee�0+i^f����[&����ݿ��wR-а���Sv�Q�룭j��������\�%1/ R�[\�ч�l���|���-��y\G�a�;t(�ۋ����j9�%�ߗ�v]l:�3+DO+U�*�%��|.��O� �+�Ѥm�,S/M�@��R�"v�Jx�I}F=y�}�%�N
<��j�䵚�p?IРʡΒ�朊�MEo�($m;2�fxc?A�y��ISK�u��/���B¹y5-�S��u���[����ôB�9���n7��z�R%Tu���*��+�s.�FU�h�3��&U0�Y�닠�Z�-�tT�]˹a
LxS�ġ�#j�2v�!G�$Xa
	b�u1zخ������u縳�$��$��@���N��«�S�=_7S��#�Q���7�H�9Wɜ&U�O�K�2��k���@L%���d�H�.�tH�l���),��epМX����+v��o�,�����4��r�ǱРCW�cf,E���Ŭ
��Z�s��:Y?�V��}Յ�!���`~ �7��za���BV�d���fިoߦyi��Q�Śo~�|OR�Z@�ns�/��iPuy�訠�ע��.�:�%�<���yJ���!��m��Y#���|%`ͦ�d
I���!��}�uG�m��wv�k�Ӹ6r���b/?��ɼgHX�$�{�f�*^��B{���2=�֨r����,m�z���a+����jh�|���Ůha5�P�E���^$2RD�{%'�'��$�GNѦ�la�8/��C� L����L�kU E��$��j����FL����[�ڱpO&�K��g���s�e��V�Λ"���Ͳ4�ڪ`�3Q�U��S��r/�[���iұ��􋑤����(;9�v�e���AJA��s��. j�"G�`� ��)J/!���0�����|&`�(&3έ�W�a��F8ƫ�B����<%Q�]:��D0D#^���q�k����V��DfJ7y,��}S�����a�Z~��-��eR����5��[sn���8/�
q��������(����	�=�6vL��ۅ*nO��R�$tGL�9P����!���Q6P1F�,CJ����?�/R$J�����_]4L��Q6����Щ�;+�|
�F�L(0�$��%���
!���m����*�6w�`x̵_vW� �Y� �4������!�ϟSf"������d�Sk�\[����y��
J�[2�Ҏ��~��E����w�T��?�}F}�@���ߡ&w�T%I$Q1�^,nC���]�jm�I�$ng��ެ ��-(��:��a�"�QO剫J9қ"T}?1�&0�	�D!ƾ�7^�AJ�᛽O}J���N	f��n-j6�����]r��U�u�����G,��v�j����5�R�ԡ�/�}����1ߝjt����>��������0g��J�ۡ�3����=dN���,-��Վ��nP�9}�h����!a�Z�,E�[�R�Z �T˜0u(ݲ$;k�V�E��Y��O4"�����ĕ ���ha,���1�����$�=*�����1��B�n����*����^+fτ���Δ�PY����a��ĊG�#��b�����1�e�.�;�a�ӜsW�8Er�&t�ԩ{��-@x�4�USl�6rp���r��Oc�pZ����ҌsJ�v�GP��[�{���'�N�-��]��-ٍ�T�'�;f��8Z�⿭�^<'���p���.��F�@����O#S3aoy�g�[o���LIU�V:��k��.� esw��b8 C�
��r^�l��N`6�C(�:=O���\�P쨼e!jm(7�^gA��Z��cA����{��|(�G�ɑs��W��.R��>���RW��r�Ç_�;�E�=~9����t�.��K�g�>Xaf�>��^��>�e�)}x߹↼�I9�6��V)l���1���w];��칭�I�?�=i"�?b4Ѧ�+S��&��`��T�M���E���^8.S�{�3;l��3UF�h�;���S �E-��Y�{Ʊ���\�$��l���m}��D
�n�G8�]���=���p�Oq��c�@�@��k�X�!�ڜ��19�-vԘi�$�N�Z;j��[+���e�9�
M�{��=�m���ie��l�E-)�����__,�^��)I7��קz�fՆ����ef�`�6/E9����4F��}�ߴ���ހ��@�O��d\��[H����r�(�p������
s����uѩS�L�llU����r^/e5lo��v��	��7��듟?}}4�Z�N��m8|i^��H�] ��E�Z�M�d_K�S�>�ߓ)QV�9[�#қI�ar�.��9��}Q1͊W_������{ ��3Z???�F��0�̩��)���&#ǜ���j��B�$�xs�X����7�L�@ΈWn��83�p���\PC;L�܆�"P*�?��п�_ܺ�!	Mo�����5��>�w��M���S�u�>E�n��~-��-���|��%�dM�4_�ܼ�hWyJ��1{:QN�;M<���>��d���G��3����=g�_W9����a�r��M_�2D�38�r�м�h Ĺ��hùv�t���EȐ[j>����+�����.��&e�\0�Wͤ�S8qc���:o}���X��B�MU�%$Ws�L/u=��ʑJ�]u�8��:�Q��M��[�:��x�,���9���>k<u���Q�E�t�/,���ip�=��NH��S���oы�M��4�R�%Ί�l�Q�/��ËP�&�?�k���"����h̾U�A"0�/.��}i;U!v�,�E�l���w8�Ν��5�)��9�R4�\:��Y�� �=�Z��u#�SJ�3�%���|ē�~�2l�8�j��:����7�`qU�O<����,�5��:��
I,޵f0���+0m_�V�s.U�-P��N?�dЦ��g�})u1~T�K�キ�ūU������W<>~�Yn��L���X�-Vz+Pf���D%����ov=��d7�9�p�K��C�3>m�3���9,��eO�\����gs�W�T�Scʑ�cX���	}|�#q��-l��ٯK��,V��in��t�5:Q��cE�es�Oh��*�ȼoSl����]�O�#�����2��ٱ=�d�NIPKY%t������O�I=���5z�i$�uQ�݋	t�_���������-��`�����٧�.�JW�p�̧^D�)���g�cq�R<x���^�7�eM�卻���V�z�"�5H~4a	
�h����r癔.�r�����J��G�|��օ�
��Q6�5��0|$�ei��5\4�1)	� \T!�4���L>_ì�Ts)}F���O�x�L�v�i����5�;��}�:�r0�P~\"�/J4VWr*�Z�����c�8��6J����*�W�����	�S�ǎ���\�����I��QU��V	��┶�Fd�����~l o6�y�d?��07��H��
M��;�fl�H�M0H �O��3�f��fm�/�������,�4� �=#BX��e��񆉂�8^ʨ�X�-+���<�%�O�T��r�c�ƫ�g��mu&��ͼ��ӱ��wn�������R{S�ڎ~�P?T�A>����B��4��J(E�w����!}�5,E}�}¯�)���_��b�����~�O�᡻r�4��ž`uk�� �g����|�	�h��+_�1�I�����]����6�_ߍ��[eݘZ�Ij�38�o��VY̦}EQq���p������&�z
�Ni�#~���@:��Z�e����3O/Y��G+&��:�����9��tq��5|:��dx��=F|�i�J6KF!0��������?�4� �`�ۜL���`�Չ�@r#��jpMl���te_�5m�*�i����oߓF�J�E�OCH���ވ��H�%қ?m�p&��j��]�CF-�L�g��V���2M���5�?y���.�"���2`s�oo�ʧaF�[�^) w
Nva��.�{S`���շ�)�`��kԸ�2ȟ��iH��u�_ׅ�ww��a	�9:����Z�m��D���|�ͩ��X�Π����6Ħ�IU���#%��ЦG^Ê��cV��M٥�yl�{үDi���N�b��rBe��a�t�[p��GQ������%J'�������=ߋ�K�y�ă�5F2���s^g�T�؎6�.7����$��sW��nw�Z���͵��Z�������R�9,�
�e]�aL��ꃧU���mɷ�=-ۨ�#ߏg�	������ܔNj�{��gM���u� }�C��O�E��j�8XC�����������F�=Vy]�9p�6yU�0���&��~��}�*�Y�Y�P 9���.M�ުrQLX'���  �i��Ok(�V9�}�+�`˰�^�@� BtF�D������$F�%4u��$���?a�fod^͋c��(�KW���	��1��C-�m�[�z�,Ƙ'W�#l�;Hl������I����!��kɯh������3 ~$���qˈYK��Z^i[��LK���m�& Ts��޽��G��-�|��Z>�]��5e�N���c�}�C��ն�e���l�P\@�Pn�a�qtO
���.�2X�95�'W)5=�O����>YirybG��v����(W=ei�w+�af��Ja��t�k��9���8�=�op���k����=U}@�tg�̸)�U�?ɜ_��,���}��-8����Q-��$|��v�\�}��Ce��)Sv��(�N����](R��Sx0o�k���;���mrp�e����YV�g�`�)z�n��}G��A^�ȴ+�8�K1����G�V��>W�P�5,�*ў���Q5��%��Y��܏Z�dϤ�������v���a�.P��B�,�]�����b��j�V�Q��v�- D��� ���H���Q���x�T����:oÔa�c�~��Q�'����g�#9�j�*�/��7�K �+�7��"������ي_!��]=�p?[5�\i��(�n��y4�̡e�.B�Iy.��w0׭C���`��k���X��i�"A𠨌�߱\�7	��:��q�8b{�ǣ���[��ы�O���~K*��h��_�m��\��C�cCvjY�L'C��D.��^]e�_������vv�%���������瘳�!��(�VK�3��ݒ�fI�~����:�X�W���˼��P�)�#r.��삎A4h�_!Xv�&@v�U^<]�ي5��e�;{|�� �?��"|+]�ɑ�ֵH��\c��;ػi�UK�S;�NMw#A%#v[� �Q����+ߗW��/i��P�-na���՝����yE@� ?(2YP'�[�������#�G��p��)�w4m6*|�I��;����";��T�dԤ,G�G:k���%��C\m�/~*�n�=�A��*Q���\�MW�7לX}��s~k%��=" �ـ^���] ���MY(h$ǉVQ���:�a���(ݙ�I��sg$X��=� 4X|�b��Bu�R~�'M�w^ü]�G�A<|�T��?��'s&�W�1�w�2��"��
�.�?�4w�igL����:�-78-~͆���xK��V݋�xȞ���ٍO1�S,��M��eC��7{�W!e����NG����׶|��_�>m��	D�Q�w�m���R�-� �����0냂��='d05	�E&��,�Y�%[dq�{�n}�	�����m�P�t��x�E���@\ٚ<��	��j��*f����!~+�1���g����>]��at��
�j�b��9�OZ����0�O�s��FSz��QʃIO�\/�a��ALk?��A�c�Ũ]���%}ld��`��x'>_�-�f��8����E\�i�ϵl�q�|r���X��|�Xq��5���#�F.�l�=�1��z�a�8Ӧ/"i[�+CA�#�����i)HX}ˑ��L(G�l�<�$y'�'���8�;���5s�C.�5��bv9̷�C�H1�,�@M��ڲ��U�̷bP�&�= �b��s�B:e�ʆ6e�-��	���b���
a3�C�)��;͎`A�O8i٨f�ae��ԝ����^M�N�o]��Gt(u=�7�������þ`��RU��q��Ł�c%��\���1�Ц~�%HM ��g�*g���z�xg�mr��(�9	�+����l�x��r����n7�A���lj�����<JXh/�^��#���d���w��aWQo���ʫ��W�)n5�C�U��e"�+�ud��W�8Wf���S�d�6?�0ߺ��
k����}�R�A�kpa!<1cI��о��T.�²ĝ��)?�߶_���~(:�ѕ���~�~��}Apʙ�+L�@��`��'�?��D�׺��qe	6	��f���?T�0���w��|%�*IN�h�J��=+�[b����2�dE�<�xʖm.F�Z1�u%�<�)�8WF����t�E��)+�o�^��]���ɐ�ʽ�L���,9ͧrp�R.��۱	�>)�NqG�Q`�s�;׸�Ad�l4x���O/2g��}�n�����Q�~�b�Ҝ���AG��"����=�&�ó=��Ӝ��ޏ�2 ⇃��6%r���և �����s�͏W�:�'N�t-m�!U��ک
�7e���&jq����נ�t�y%�JDZ�u�IdJW�S����w:Z�q�|]6���˷~2��K�+��w ��;#��8���|6q>w348��i˚���J���4A�P~p� w����5���H�Y���Pa�b��O���s�t�8Ӣ��u<H�a����;\�Fb�`],����-呼�&&� �nn9 ���*�9^1��4i&�Vn�NԪ*p����(c#��/��H~��$������W�H������:�uP8K��ڂ/�"uA'�B��[b#	F����pA|����c�L�j@+�ăxL�8If�<�%���X<b+��5}w��^�̓{�CvhG	��^_Q�5lݟ^��Z4[�#��0�!��!����W)�B�:5a,!i�q��Y�x�}������V2r�Sh�;����jdZ�z��}L�8Ο$�UH�ͼ�>�T�Рtٹ���������\�F:�}>�����.PX�U-�Ī�A`֖n��_`m�S�pO��В��ڠ���L���D��.)���Y/�V�R�-�b�U�L�uf�Z۟U�v�rr�.;S�|Y��	eЧR�ѭ<�0�
�LK2r`���T��uih��j��N�o�{�x�G����4�^H��$�K<fX�׬���ɬ��u<^7�Ġ14��+Q_FJb[:�;�eя�2wI"[�I�AW������bf]���/���/כ�Y���Ê��8[2����
��Q��>pA���
z*i���k��6�V�!Ħc"�����4b�o����8O�V0���ξ� u/��|�,��/,e)�5�zQ����d�!k�̮ʣ�i,
a����;��³v��X���nHF�"c�ر��F&.ڷb�]<�6��B�@v�ۚ{�3d*�5��
�g��.����iD�fM@���튩�{��<{+L�����ܝ
�G����Y��?|��k7�`5���꟠!N`��t��Y ���d����R5XW*/UzI9>}� ������ )�S1{=�}:|&R-��ӆ�^��4���R?�sz�2���g7l�t�����.^t]���F�<Pi;�QqF�6�},�Dz��B�M�e���=�3>�ȗJ+�I���Z��_����(��e ��\��H��Q��F�xp�=l������x�.����)&�� �?]/�o�����_�b5C��Z)^��\��~M�s���`Z)i�7����<�����w��Er��.��U��J�[IA'O@X~^��w�@�`�KǙ'������M鄻�W��KaX�R�[�Ϲ�5��^TѲ�j����Gb�f"�1H�W.ٙ(��_� �]d��G8�M�N�[(�i,��8�@����fDe\�������/E�s`��?򁊜�q��'����gErPr���*���J�w�d� ' ��W�_�R��zc�i����j��g�o"ĺ�^4��W��Ȧ�Q�J8!)����]p�V���	�qL�w���W�@��g{X�v�����P%�:$�\�����I��o%�suxO��-hٻF�X��;�]�� �O��N�|�Dz��]�"�HC�l�~�/���Q���`"�l���GwdIb�Q,Lu�$�<�~$\�}���X-�(9�ܸ�ǯ4wy,��Vo�����4�g�r��?}�j���{�kU������@�R��Dќ٠۳7^�eӳA܃�G2���qZi�^[@��c�rY8{q��`�>��JD��������)#�L�s��~��H)C�u͜=J�xHRE��z�m*ݓ�C^�&k���u	j�����fe)A�h���M&ECd
�eR܀����H�0qI>�(<������_��G[���9��+q�#L7�L���:���l�0���D�7�!y�:������ Óf U��H�L�s&u��*)��v0��u��"���4�:bI���5�n�~x�#Moh��:�e��,q�WĒ��s��,�6����C����P�7�Q'cƑ��RP���ro�����gW�'Qv�:N�j���`B��D���f>���u�ؒv���n�Pņv�z������dC�� ̙e�qC:~ޮ�wd���2���~i}$��ބC�&��s��gG���{�%�=V��kd�{��J�T`�CIK�S$�s�v�Q|ͤ4z ͇��m�����`iV�vR��4\+�B��Z�{TQp�w���t�MSm[r�}-��V���?t����;^a1�z��
��#M�k>!�OY�#yݞ��Q�q��c:�������e��d{��+\�%��0S$=%�2�2-������`�<��8�'\f��` ��o�W$s���k����|��m�����Kx�$��:�g��җ�LvPZ�'R����R�p���Md某s�m���\C�黚�Θy}��0����7ڤ�KrΗ'���.���pY�N�B���B2 �WO�}�ڞ2��~��g�dH]�},�Z����v"�i��`���}��E6��?r-�y�s�'��+˸���MI�_~���rB7�5�½MT�;�6��d���*�� ���2�Õ��Ũ��%��L2#�e]�E�L�/$:d/F�EN�e��.�?�S�hRѩ��"�pB^�=��ژ�Ѹ�X�/"w��ؚO�qw�4��&j�f7���?��C�>�A��u�H�>_��`�$�WSkᬱ���
h��e�ȵa�䗶�t�,����Z@m��C���4��R���<��8��
�����Rk
Zj9+2�L�c_�!�^O?�T�q��f��E��C۹��GU��UH�$Mu%[����YQ:��W~[ษ-�-I�#�&���᮵H�1�������Fi�Ԟ��n(��_�;`UN��u^�4��;�]ؐk[gO�g�t�6Ș�����u�Z4B�F-緕L��A�%&���p캪�nSWշ�\�e4n�`i��'U]��y>(!{~ '�(�`�x�ȥ6��CZ�/!���ju�뎨ϱϦ�����GGA�_�%��J	���8�_�uq&�W�Q�I��N�\d�z���<��DW[|�
���>~!c�Y@�j�#�7	3X0&�����R5�R���}���y�y��q�r�|[�T;��_���@*+e���y�Zy��._�W��V��`@D�D���ĩ�4���ӃO�o�IK�	��R"��켡�(*�N�������Ŭ��U���Ԅv��@Y�%�s@b�]K@�.
H���.��w�oV��|"pe!��=�H��X�U�<���m���?�Y!c!���$���P�t���sA�߁�Z��}i`X9L�+ k�ݥT3EX	���A �Ȟ�i�W��_���%��[sY���?3�KZ�2T�[�h���9���~ox�����W�3!2�b`��HQnH�)/g{0k8�o�&���+X�J;m�R��D�YfF�!:ј�i
�k�.䴢H:�
�Gu)�#(��2�/G�6;O0����%}&�i3�z�?��RN��H�^V�����D��VI��}讫�!�[e�v����r�����)�3���L��z���8��� 󌐾�pI�}�mzJ���-��x��P�<�On��:�ȕ[?S���"z������ڞ툂�4t���҃CFE�z_u6�mO9V��ΰ��5��[��#��e���uЯ���]Vʏ���L�h�/����C�}t0J��'��~^v(��n�2��iY^>���?��:�h3r^.��������[����8�^l�-dݪ�#5��@@����P��@��&�I��Ot,JT�� ���-2Ua5��,i�� 8_�`��,[n���yc��G�΍pO�d�R����ƵSs��w�W��@&o:�ťE&��ά��q�&=-O��5KP[��E�hc���h���4E�i�~��ͼ�y�d�w�e�ln���?�uY�~E�	�$^1b{�Iy����:���Q�n���չ�"u���'���hK��չ�T�kt��EqXL%�)RU]9ܦ�>�w��SA�\1P��:��	Pܪ�/��ˡ7A�w�����=C�U�膺�;9�}h�cC��/<Ċ�{n��	��ǚLP.��w�����OH~m" ��eBh��*��_+I�By�3��'W!�=��� d�&�2���Q �LW��R{?r8W�~iշ�Oƴ�*]�1��ǐTT܀�D�P��`��t����5�
$�DOI]/�X�V�K� t���pt1����#U�~�f���-�?���#�t�]�����~B7�8~�1�N��u��NISJu� ��@�X�e���:L�uX�k�"?�o�AS�	�ɷ�{�"��x��49paǉù��)H]�Q&'׵vбk�E���2jBo��x��D�d�>�(���<��kX;���!�Ȼ�$�~[?��j��F�yw!n�]�x����aW��h=E�U��4�*[����Y%BB�I�4�U��Ϙ`�;���Ϩ�a�:�h�7��C��5��e.���9�0M� b��e��C��i����.;��DY�=���%3�%�"����z]td:�E����3]5C"Y��qիP+�<^-4?\R�x'WE[k���4��5�s��mÍ8t��"t�@�`�P�,�桖� N����Y}�-[��&�F�Ty6�Tw�97��s��;ɖ?hH&���'4���h�Sy����F������`p&����P���\�.䷑��>����b��X��i�K�>�n�#�Lb�,4Dh�i�c7�Ƃ	;�̊4'@�����_>���*�sύ?Io��7��� ?�1)�8@M�q���?�n��ero�Ʈ'�%,b�G�g��n�g�x�D���Xd%*����n��1}�~�,w~�ԡ�f-��˭x/��	��j��nN���e�Z�K����H*9��b,eo�Rߍz����9W"0�������������Q����:�Pj냨pצ�%(���x�%���.}o7�m��o(o2�Z(�FS�����9��$��}�������o�&�E��-�h�Ԧ���J
��6�њ;���/���82��mm�beik��t����p;���j���h8Fk8u4�HDog&z\��o�˟���0e��T��ћ��g�Y[�+�}L�uO�RR;9^4�#�:V�,�qLq

�l<�l�󘞻 h=�5�U�$D��dGa�9S���u[S�g�&�&�
D��A�l��{b���ёyL��
�3��K��rF�X���/\�G�� P��ؒgn�R�X��[<�3U�#n�.�6t���v}S��r�*~� z��B���M\+/V*�~n,X���_�����
+�5��y�)a�V�آ��R	`�:,rv:,-��6op��~��0%{f�G�>(��#�0�=&8�z�-e~S�����||M�H�\�r��"����a�ٔzʞ�Z�m��.B���{gԍ�WV�rd��Lg'�띿���=����(�����d�<-�2�6��zKv�r���`p#/���i1h�!V������;YR�4鴑�{�&���z�K)/¥�ޡ� ����E�cJ@,�*��/cz5q@�:��'�H�"�)Y?K'������� 燎�W�C��UQ���	���rv��3�Nn$�r�@;}Л���GL���}�����#�*��X�%���M�c~�7�cu}��S�y3�h��r�\2n��T�xy�v̖P%��|���٩1���0Ȫ&d�L9���Y�v�ﲎ|�����-Φ��E��@:B���[�B�B���*�}��슢qow����l���?��xf�g!�)��auEv;�y(y�GB��c?������u�-�8H*_���R�bv��� _�lw�m$C��gy�z����٫�ߍ�E�K� �	lW�κP�@˿��W�8|!w3�	�t�O���3E�%4��JE�N��>���n*��&6�q�+����1s��x��RU�˳KV(���m�a�Ű*�z�+�~�����T����Nc�l\ �=MJNkр�����:õ��J#Sy8^
q#7pT���w.(���Z?q���;�L� �h^�|��{��u®I�	�>�lK���]F�S�Ih�L��}�Q54�Z�@�nwjk~)�Tx2:{n��`��l#�+�����@w�y�7�Qj��P�C��w�xDiӁMm�uv�n����а��H����*���ģ�
K��:5�<.�x� Q�������h�NJ���_c�8�B�T�b��J�ف���|P��*�r�D�)v�]�����^�o���A��2�G_��r������MɠF�>WC*I�'S6�|����z>f,�!�N���x6�<?�R��r4	����SL7z�����$d5�\�]�%3��V�n���[��>���f@| ��V�Y;����S<���{����&�l��e��D�/L�E�?b�Ǡ�G-����K���bT�k<o�3�}ŷ���moH�]���:���'Bv�D�V:��PE���vKB�h>0������sɀg�W&�@s$��HM>�Rv&\����Gxl���)&2�k�.���Z� Иa9�=���+쌜�����c%����7��8w��~����3:���my~x���4�:K�3|nu#��b�T)ܯA���7�z�z��u��'�$�=�1���;�i'��".2B-R�ÝDD ��~���F�O���x��w��f=�����e�ė�^j��[�!pB�EKr읹$Bz��F/�~��ϔv��Nxc�Ž���5���_D��]u���}q��E�ҝ*:�`�|~�� 4Oַ����7�I�����L��c��k����;ițyi�Bڙ�B�l�=w�b����FH�p�m=*:���yo���7��(�&%>'�]�\�w@���	WU��\D5�v�P@����a*uēaH�&��Z������H�C��D(�3cT���5���+)�W��Ee��k���1~���DT����e�j(c1
����(�yv��qx�@��TWS0��+pmm)��k�k}����t�W�P��ëM�L��J���m��T.U_�+�{���TgYpLz��c"޷/
�ou����[8BAa��;:+��'@�����x�Ҋ�fc��q%ʠZ�&�����4��������3 �N9��܈&zğ�e�C����-}����i���ȷ�yj�B�r⼃�$l�ɍչ5�cM��O�Ao�(�%�>B��m\����@-��g��tE���sY�^y�k�H(7�����1G�=�r]w�y��C�0Nl^V�y�Wf���v�i�zR�#3R����0�TvX3V��ՓCR�N���Lc�A�sy�`�r���J�"�N�kA�:n�]*�'o�1��(�~�<]�W��?B�X!��Q�)��s" 5�+��.T椕r��@��a��a5�W@��L�^;è��Peʪ}.S3	��%�x���qg�V{��\Y���=]�&%C���
�nd������J���ϵ��>�2R���-�W�Q �e%��~I��0�kL��Ir�RXْ���Q4?�v��G*O���<*L+�.�?�K'	=�SH�	H
��#�,���Z6 �����i�^>�׳xl�Oc�H�~2|J_���ʧm���=�KU�2������q�g+-�a���p\OPb����3�*[�r�]	@��!ey!����x����dg��i�<�����H�(�*��������u��3�ѝ�ωj1���~���zY��3��~�eҾ�	�YN&�f9�DШ��#T��+�����P�#��4֤���ʜJ5B��?i��(�R����6
�u����wv{����
�u�9�B�V���:�|���}�^�#��f�LڌS%˾dX�X �b�x�]$�MV����~�M�4O|��{ �os���༦��O��S��k��
��U�&�����4�
�hND�4d������L޼":�-8m�Ŭ�Y)�7J�z}Rŷ��[�xKN����UkL�`�bzג�":�!��!,�7f��V}:�����'q�@Y]������~�̓xw�_� c���.�a�p̬�h݊�^e�x�XF��Zm_�TA�M��uL�V��(�8�?��p͊�Չ%��M҃����x}�G�X�+u���h�^,g���m�P�����+7:;��a��+�@�S��A6)rĬU���f�
�e��̖O����گ��/+���)��������֡�Z��K6{/�7U��7���g@v���e� 	��zH�6�����&����6���ߗ�yZ�I���L.���w�U�pY(`2샅J"�'8&�m�Z	��t2d�x9��R|y�+�S�V�-���%�7��,�K��$�����U�c
�Ƽ�p3����ts�.s +�b�^
���J-������09�rE���S����,<3>GtzO�)~�k�Ѫ�r��	�5��-��9p�ڟ@cx�F�����"�(��}��*C�qI	�c�m[kc���}�.蜚���ь���aZ��T����+��	FFH4���hC����������?��|Z���Z�#�y��ъ�����3[�D�o_� )�1���/���sv0p?R��p���6� tL�`mW�k��N��k�y�����ׂ4JM������3l[)���l��Uc\�s������P��_�6xKW</�X���M��yR�81_�k/G�V);�q���3�&��d%�ޚ汖���b��5�7�zxz�<s�������q�s�b��91ƫ���;o��nh��T~��L�5[l�
(S~���	V�"���$˪?���^}�>f�ăq	֎O5=+1��0q��sF���(��ͮggUg{%���젎u5ʠ�h�%�2�P�h��3�:󻁩X����EI�.�s�T�bO�ee���HE�>g-����OXc�8�vf%�`��TDiu�t�c�v������R'Q�����#|�#dRL����֖�pE���F�������i<y���39��h_	��	$�^d�o9����&�ڕE�����N�o�����cmRF�g`,��+i'W�{#K kB�-s&q�)�CPī1[w�'(�Pi� ����E���?��@+~�W(���7���Z4�,��xK(��~��Ʊ"k��T��]ٮ��$��]s)�ե׫[K����^��<�ҏ751���<@)��*Q���r�*�6��u�d��@�e��Hh�Y�j�$�r�k604�2�y�zo�����G�|��� L�f�ۥ���A}�e��n��
�#1ڤ/����E��sº>F�v��1-(�6���h���J����Y����c�@Z�hK�E�ھLZ�_��
�SPՃ���u�}`]"Vɞiq"���C?����F�0��kA�,�{��<�32\�Z*+/��?�;�7�����3����P����I�]��^B��^���ޑ����^���i\��_��p�^ү#19:�H�՚�'0JO�ir�FBN�Ѫ�	��7kj]�H���,����홖��̺s&�cajpkO{���p�[�zlx���zט�#%�R �?@�����i:���Jz�e�8��,��
��(G���l�y$
�D����ǁ���gzf�I�q�C��L��a�ɾ''L�Z��,z�i��\���;F$7].��Z�6N��on?2 h\�k�ȣ1��=^^�T��ݓ�h��2�^I���6_L>��v�r��i�F�A���I���-�h橑�hշ�5��s9,�����E�pV�^�)��R	�d�V[�^Tļ
Q�uk*��x��k�/����IAC8�?ђ޻�K�T��sxm�-q*D�"H{Waq\��8i���}�N�8�X��p�'/�XzX*��M�aQ�)�.�Z�"+0��ȱ�)�mQJ�2�(�4���x��([i�����'�~C���x����t�C��b�f�lѤ:{[��<�([UL�[�|��a<�3��+����:?��?W��?�W��`�r���C��}�b�/��szIi~2V����Y;����j�q#������:�ƚ�\]"����Fk�k��4t�RQ*�j�S�ϛ�@-=���Hz7����Q�F��!i+jc-:���үt/��g���C����l��-�3X������&P���.�π���VmM�k�8�O�
xg����<x��A�@�����0s�=+yJ�2���Գ�� Dq�q��$��e[����$)4�G�����yt�Ɏ��L"L���|����9��I��kԡ��>{I4�bU�W�p�,���n��K� |�z��t����Śı���eE�%��#���Tz�K��:M��M��~���/ȐE�,���0գ3�]p*6�����#,Ngt^�"8�Xs���v�v��叙I;��uR�Yz��aI�C��co���Fӟ�(9}��I\ϡ�JB��9i��{��C0#k�������#s��3pۘFc&t���e]*eyrk�_mo�h�n����4��ҏj+�2�KL�$�[|��p���w�Q0�ڭ8Q(����+�p. �㮿o�;�p��줅��P���dqH}�z���+�sn�㝇2G�P5T#4�kؓ8fB��bi��G��e0Ce��D4���	���b�_4�>i�#�#@�bL'Mr�⚲_wZjR��O�Q�I������}XW�gW��5t��%f
7xF� ��+�w|�m~�6�U�cQ�/<�D�2=z�қtr�\/��aZ��g��wM�,��<V�"�hA	J��ߚ�i��j{�̣�}ߵ3
f�`����vȭ��;#)$�*�
�\�,cKT�%�Q(g9���d�f�#�-���C4�'|���5ֽډ��n�]:o	�(�.����,��߲��L$���i���rJ-��e������a��b�W��b�i���)����YR�����0�*9>r�ݣ��`�V%]V�刺�����ǥ����l�8!Y�/�St����&�����P���$�����|Rd�Mt�:(�_b�#�OЪ�m��W'I��T\mf��BE� ��tS"����{�x�P�=ř:jv�j�'ˏ�ŖL�ٯ���e�Ș<�x��M>��5e���f�B���FuC�����mү롚������Y�ٰuU	n�)�����e}�?��|����N�!�EA�5?!V�0u:���T�Mצ4�HU�}�gCjm�G�՘��v�uc������(����t��͐��J&?�ܜc=@ip*�_T���Va}FpZ�r�UI�q��ۗ�3�u�"r�v��(-�|n�!�=�������#d�9�GA�/�S�4�~�W�q��:}ε��k��'!뮕�7�=��9d���Ԝ�ٳ�P_��C�WQ����T���5�8�V�k�S?��Yi�4(!�}�8G�CrC�s�L��3������-���t�y$7�)@�^��U��Ő�4�ˬ�8�9�`���N7�����K�_������A���0��0���r�ԅ���D$�u]�w���n�N�szs��I�R�;�L�j�\�̏��֣p���z"*0�ƒ���������a:�K\m�m�gi����Ӡ��<π���X����^]�F��x�2;e�3L>x�X��M�E���z:g�jL�b�,x��9b����ݴwKr�b�I<��E �+y*<�a���x��Iͯ���z��5俷B�O�\=<$�8�L	���x�}q��i������4�e!�9~t������[�}�
<ob0UԲ������R�B��/��x�(+a�ll��V�/˽�>��9�}$%(S��Ѵ�N��zaCZ�N��]ߐ���dH������ A5��p ���Uϯ�nm�K�>�R��{�8��>�O�����**����c?���ׅ��ǺH�X��N(dᰣ`��95����	A�N8v�us�s��G�a>j�Ϣɩ����9���+���K��?� �4Xj�db����kw�8���0+��Y��۹�
�
Eϩ��d�H��_J������5���cY����;�_�.�g;�Ӫ ����*j�[D|k6���񯜔Z{�x��`�;	��J�DU=��#������ �������1+=��%��G�����[9Kc֮�f�'˽jE��?�M�h����>���q�"�!I�×:�B�ʍQ¦_`�s2�*Ģ�)�J�U��i�ߊym��/� 	��֌LH]}b��,ˉ��wZ�gG�[�o� ��l��]�������M��x!�FF3@�֡t�8�cҐ&�&�G������w�QA��:v]�L��;&W�=�t`h8��)��6l�3����u�0�Z�O���~4<nYh~�Y��O��Q�LE'��Ʒ�1���_����ϊ�b��#t������_�H�������a�1J�A6<i��Q*�� /�:Ac�wv���>���sVrxo_V��d"ጰ��e�A���h�i٨_ǋ�]n��ƺ7N�ؙ� o�8��n�:�S�t`�i�UX]å�)9�ڭ~��:�
l�%��Pn�P��ps��W~!P�v�!��I���9���䤬(�Ѹ��E��J�0XH�y��<����qll_����!�2�47P�ѬJ�:+���3�pʁ­�)�c"�l���SGCJ�ifM1�����̃0m���b�{���R[����#`E��t����Vۙ��4�ˡ�3N%η|	n�h���,��ԭ�j3���E��Vo� `L��<�ڀL���ys�	iO���ڼER�{� +-"8�AL��}XJy�W#�Mv׾ZY��f}����@\����o9I�<�'�/��!��De������έ�y�s�
t�9�{���O��&��m	h}$j�;'o�����Ɩ���8���!�q��v�ZO�0s}������B�oWN<nN��g ��*w6<��Tp��S���,� qF`�Y�ӳ_	�GNlؿ�� ���F�q�ߝq�<$�%bw����fs�WO1�%�=��2��?]�vz3=�W�#�ݤy��m��ϻ��1��d��M���58f�{��d�ԘoS�Y�F��3�´�>�,\���~�2O�e;�m�]|��o�9s%���NV)��L����Ƒ�uh˛^O��i���u���!,a��ہ�֜a~{�a�q\
��@���8��T(UBn��x��tz� cU\43��?�_�iƁZ�ny`5�@MJT*��F�������4���m�m[��惏���o"�q�^�� �z���]͓w�,����P�fޡ�f�ߚ�)f(c�G�vxh)PY�ea{�]��G,8 ��]��?�/�t����{�͵���VFl!���_%m���M�kM�dIz܏;U4h����!E��;�%��*��� �b����H��~�<��܅�ϥo\��,���1��X~�3�\�os�w��+�bM�C�<���x��@�A��W�����(A�9��KB�g��`�x'3\z+�y�(�(�N� }c�uK����*�<:;=��ĖI���l�U�4t[SF��0DΖ;�<f/�wz���F��Gvu��/8.��#0I�)0�ʜ�œ� Y$:��:V�ɒ���;j�iNj����7<�Qu�8d����v�8�a�Y1�g���r#�	����bZ�d�����P�X%��ݶ�\d����yO�5�ӖC/r�v��Z7�$� �Q�Ѿa!�����EenhM#m�����>�	�Ǉ�8 �` `�f+�I�4H>�tr���{4�0!���C_�rj�V4Y[:(�vyhU�k�(���>8���bJ�6����-��5D�1LX�F�"�Ī|g�U�I��d�|��Y�r���k��5����JJ`q���4��"tѧ�w �J�y���-o*����匆jޱ�[�0w��?`t���26��^�(8s��n�`�=�A�OfX�ͨ���8ݥ�ˆ^��@Ѧ�B�߬�d��(Ye=���_�F6w��4h��b?p��tb2H�ZX���;��B�>�"�<M�}��ȑ���9�=�{�s�SX�~P��/xe�����x/Up/���ۚY�7p�zV���7�����^�^��v��ԡ�)�@hP��.O��p��O�3���������&$�:�f���Ӣ��z���M�R�gڃ�ԟ��o�sִH�fM�r���H��}PD���>j&A�¤ �_� %��:��͖�����y)V��f`#�u��cf��abB����L��F�$��sm��S`��Gk�T�M2��Y��G|�X[yCq��i���/'������j����l����u�4�v"8����3���EOٜQ�^kH��W�n�)F}�P��_LD���#�dA̕��Xp�`�۰���<x�"[�)V��P��r�.`>�]�#3��w����H�鮶�N!�'?�f���sP�#�΁th�T�u��u��G��~S]ui�Z!2ڦO`�H��r�>i�����f���i�Y��Kl���z>*��Z��K:k���cϮ��XJ�=P1(a��b׭8*�C��'���Gu�:�[����rQ�T��±֌��f`N�wC��LKm��E59� �t^d�����w�����9�f?�JƄ��lHJd�Vy)��CTS��L�=X�4/"R˶����n��k��h����s�O���hʞ�M�8��lq9K�EIg�� ��bm�ރ��h��f�A`��F���>�^���ɩ�p&�R�:�ONU�� ��`�<o�`�wM��KoI̩ ��I.�����k��eײ
�>f�~A�*��)����-�h+C�V�*�4.u��!E� G�jD�Y}OԘ��y5��r8�E�b��;�.�8�B�bvsz�
��E�cBt9F������hR������n�j�S&5��x�=�T�O�E=4�^�CZ+5	����8���чs_*_X�4#T(j!�,"ɉ6�eS���R�|V�̽HB�}�L�b�c�D����j���bb���I+��wr�گ��h-�K0���|4� 0�p�6~�Z�NZ�n� `m$X����K���u�����Ɋ6'LrFP1͋t!�a��\�AK���B����A�����ex7�H���J���8�]���f�l��5��{���9���zX���=���sx�3I1B�Ρ�A�ޕ}5i�ݐ���y@������ �.r]��������%VX�u��~X�aN|aȗv*��/�ÇܵC8��_I�EO���f�"T>���=��p>���+%�\�fI{����,#���ڌ��W�9�k��ڊ$��^53l�����r��A�-tD�N'4�,���獌�sA:�V���7k��7n�Y�M�T�Q��x���}(�Ɨ=����f�1�7_�e�-�l�8w�Z"�z<y��	�FA���չ�U�P��Z�F:J���B��-/%��7:�-|�w��u����v3%���Z��ȯ~BZ��dm_�|q#	�<�h�5byʗ;Z��}�?u�>��뻶�͈H��V"N/)��4�w��@�e��+��F��37��&4]X�3w�Q �f�埀 �����9��pE,̓~�-��z6���vɨ�bBa��ׇJi�0�{�h�L�T�Ǎ"[6@���9�<k�!�t�S����4��+n��`��'ڑ08H/nm�TZ���q�'���F��!SĈ	�!tcĈm�~H<s��/���Xl���s8GgW����V�6x��Fd��D:�<�/,lɈ���ɂ�eMc�h�N�%Q_&��W�i�;�'K���[77����+>��	K��K�j�k�@�{�Tw�f���_�d-�M5TPb�������H��_�k�Ϭ}�����(gN�'S�;�/��Eg�t8x�z�7�����x���P�"��z<�J��s�;���C����6�0�����FUЧ���a�}�����\\>�P�(�,�h׉Y�����������fF��C�<�ɜ��z)��r0g���#�DO�X���J��'$*%`��:0�k�X
�lb@�+��G�KZϘeNbf쥘^!��l	�&��\KxPe���Z=�7	3厱�_���mIm�z�L�.��i��"�I%���|�δ�7�T�D	1�}\�S��F��fJ�=��7: ���,[M��n:3F0�p��'�����B���8V�}�mzO�|T�/WV��v��"�v T�9 ���z
IJ6�c�k�\U��+C��$?[��>�:~U��+2�ޘ���З��x���H�ĉ0�*B{���4`m?�*:��C*a��]��ɀ�`�ޕ7]���y��OG��7\3�c���;0��Vh���TO ��#�$�vk3��u&�o�Or83��T�VhF3��*{O�s���X���������t �YN��*^]�(���� �V.��f�mz]�*��]��a!�5�^J�h�v�	dV�(��h�H���X���c3��<Y􏞩��3�� m�W�O
�(�D� qϭ:�K./�7�P�;>�.�th��$��/z'ڨ���{���0p{���\�����Z<���-��RPJH��pB��`�F��7�p>�g?4�L�6R�gs���9�di�#질��e���Tt�� 3�8�D�i�-Lc�o����[��Ww����=�O����E�S����t��0�W&;��&GjCQ5՝D�;kA�k��8�9w��H��bR"}i����=dn�v8BN�ѫ�����F���	�x�F��e��]VC�7����P���qmUi�^��.A<����@)ԍbWI�ǚ�e�-n3/�Hx��T9"�H�>�{��k�Y��ty_�9����8�k���V���/I��(B1��&���WlPG���-���W��Z��Y*/�P����`+e]�3���Ӎ���Ф�� é��_&�l�����)��K�x��DY��9�;YM֣X���ϑC�����Jh?�Jج��-�v��P��S����h$ٞu�)��8<}�;;W+4�-����yc�1�O�uo��U/�I����U<9�(�ύu	L3w���9�Ұ��ꗌ��n�94?4`Jnj����V9r�T���E�)d��l湺�$Sy�J4'������&1w���潓���B.N������#���|�fP�� Mb�|(�>ܷ�t�(H$��n����?����W�(����-����D*�k��=LsF�i��n�{�>����mW���"�X�L&����1z�q7΀L�$���G�Ѯ#|�"5L�y�R�:f���`�qK�3��֭<���8���<�@0�'�����] ��B��@{�3ʜط�j'�	�S��P��l��� ��A�X��?=��b@<ސ���]؃�^�P��"����hQ���0�[�}`2�d��v�� �	���U�2�5��;��3]*zWiI8������e�#	����"�#y ��0D��B�,C=v�[5����Gݙ�H���N���)��d��w2^�Z��A	3^�H��Ն�����,���k�k�/�/S��I�����]Nu٥� �S7��8�l�:�o*w#7'�dH�����!�b6l�%���^��/?"ZzNR��`\C��/�|��@uś��H`��������*	xlR@�é�C<fn�SPJ9�R�w��͊yqW�����6��	BV�WgӴ�Y�#�`s�*�l3^�!����1�r�Y}O�m���j��d���VS��i��v�sd�� lГ<Y�,���L {�<��]eIXMS/��.J�p�&t?���aL��-��稀$�G6[?`�G0Joh~�o���ۏ[���N^��6���;�ڢ�.ox\��~:�zZ?�:�/��;���*� �w�V�m�Tj}��`ǥ@��YC�<�C81Hh�#zY-�[���-b0������b��r;�S�����l�P�4o�}�s�j�i�^~z�h�bXeh�	3�[�����af|���\���Tʣ�ao���u߻�Ɵke�G��x�O���;L��F������y���'��w�ݘ6�/����x�JF?3�s|�Ѻ��!�R�Mj���#�J�e�u��cЛjH�Ȑ��*9OY�:t�[H!&n�����t�IK��+Z�X�}��Ei7l+�I��ú��Q�����n�s�	�}#���\�	��<o�(r4T ��x��n�d%�i00��������ߞftf�8���f�b�U����^�5/�
�A�qP��(#���H�%�y��Kg[��6��.�.I�K�������8���{�|�.��gW�p��r��CH�s�E��K@%vRP��S,g�K2��Mt�_�8����Hgƙ��[�������v�{j�/��i�w��C�P��HQ�����	��uC���c�8 ��.�?��3^1A���ɤ	O�󲈀wd��i�X�X�t��qHyl��uwRrP��r�˒�ԋ���;D�k#F���3H��H���x�
ʵ��\��C@�|<�!��ŝ�Uׁ�bnb$���k���J�Al���']�]��^�?�I����ȵ���M%��8���_���[2:_�a���/l.P���x}��8��w��60y2��(�G��
O[�֑��ʗ�9}������_�J���k�����?~��g�e���kv��0��ck\3�MO�#���T��?}x{H##�廆�o��_�S�ߺJ~��o�cw�Gf�}_0�������z#ǝn�D�㜯�T���I�����c��Ԓo�19��r��[�F���K��h#��<���f��L�m7ͧ�p����G��劷����آ.��t�t�Rk�B�/��F��4�����q�=�F�رn��<�j
��3������8XD���2�ٔ�@Z�x/�k�<���Qg0�{�<0��,�t|� �e����/e5��9��E7S���e����t���jC[�M+=��}F l"�C���7>|�0l����b�ƌ�`���F�p���	�Tw~��yhhJUL�`��]�g���xM�a��@A�:.�]B^"E���fU�:go���2aJ�]�a�yn$�o~��.U�5T��Վ{�A)�M�9`�	��p|3�n�4.���"�>Ot<�,�73��z�1��n�(z�%v��lNe7.�L��A��\���J��V�Ε��c��aOz-{L�|)��?d�K���գ�����G�f�����!fK����+��R��8O�G�`�/�<�l�4�%?�c��ѡ��<pS���21b��,�)E��5�3&�$է9�Q���%Q��Δ(��	�
u�����7
�0:��-�m���x�p�l��6���~�?��Wëꨛ��~�ȷ�R����2Y�%��ǽ�ՁP-HI�{Q��#�鉢d��#�y�Y���T�W�0�ŗ�{�c��V�r��P�c�N��tT����.���c�P~t:�[_ɰ���&���r=�V(�)�>�Z�S�\B){�v�d����[H����3+��/���Vdp��)�	|�	iqwk�#��Wǘ�O���U�p /k��1��"ZMHJimAxZ������64�$��X�c��i���nugo H�k��Q��0y�8NRv$ӓ���L��6���Ze.`�u
u�9g��՟cD�ړU�}�̩����ʎ'�lh��� Zqw����"���b�=y{�x�Y�gd��+��]w�P�w��*�Cm��$)U\9�س����ɶ/������ӔY��]\���c�2q�XZhf����� @b�v�^���f���[b��1h;+$��鋾)�*g�ds��������������`H���+��I��M��A���i�:�|N�C^��K!�8J>�쉩����n��_G��,�F�f���6���:
�-��*�9:]	O���A9P��X*hص@9EA�����+l��嫻=�ݔ���/��� 3�Y���kq\�Q��l��w��}�	���\��.[Ҝ�W�}�@N�'���z���Y'p���~T5�݌�Ek[����Y@?�rl�t���B�xD\��n*��\�leK���-|���9��W���b����
������"��Ê��6L�����Y�1G�ތ�Q����P���\�̸:D���Cj����*�.��B��a��Sz�f� �"�^{�>�D�� L���������q6�*5�1	N��8�7%�\��ax��0��#Zr�Rg)*ƱwWg��ٽD�y5�$c�a�9w��Z������L��_�"�X�'hp�ח����[�ђ'&�Q%z8 ^�(EJn��[�1/f�%=�QEM�v)��?~@�b��'|��w��Ұ/�q�)2R��!�a~�|.2S�4͙@����o�Psk�c>��P�`��R���I��+������y��%+���vQ�'{�ml�E~N�=a�N��敡�:�OӜ-��9�F���1�G���ҁe��^8��@�`���
��Vٜ�O�k�kBT��F) q��Y1���oic������u��c�!7b*���3��Pe�(�J>� ��.����V"����V�^�n��g��̅�m���9�:, 49��Cp+g��E
F~+�Fyڧɐ4��7}�w�;TC�p��R����t9*z� ԭJ�7��)��Za�����!{ʭ'��?��
���?|�||����<�`bfm|l�%O)s�߇����US��1������W����yۃ3_���'ã.�+��U���r�Bt�հ=I���e�T ��OC{�qo$�Ê���>X�S�#Īp}��WY�%����a��d�}=bf/�ҜF��j��+s=1p�3�O���\�XC�'�����yU�"|�8�uQ��)���^��!��i��N��a���P?lusby�&����\;��!w�g1,_��k���U׽4��(�ˮ�rθL��
�g� ��;��.n;���%u;IMQ��-�wB�0�?�k�΃�F�_hś6�����%�z��2�G�x0H�`��/��C���La��iY��@����������:C派�D�s��I����n��&�G�Q+;����W�f��2ӯ�o&H[e�ȿbå� ��T�:H����/i�J�_�<�٧����̟��ls;a\#ʏi}�r�����C%팽��t�;2�1�2�}��F�@��A��R|Y�Ǻ���������g��"ŗ�Ѻ��Z�Ř���ٶ�b�κq�����&t��P���c��ָPxN."���N��#OcV;U��#ő�������Kؤ�iRT���1�\a���>�;�r?c�#2����>A�6��w�����#�z��Ev�Z��ӰZ�':��'� �����T�rÏv:��k")�'\��
m���_v��$ƞ�MVR�Y���!mc	�U��e=��o�ޓ����_J��g�� ��\�p�r�zn�m�IF���{���3��wGնdc^�2����E�OܼQ<��p�˗�lp���f��߆O�l���:��(,��s�04��}��BwB0���|�p;e���B��s0�Z�q���?�h.N�����4xG���d�����I��]%AZ����O��[5�o����y��IBe'ˎ'�Y�:��H�IP����A�֦%�Ũ*�(�h��o+
�e��C���;�J74�9
�>��Wh�+�cV�T/�J��3j��#g�@Pgp��^���~<�9��e��|Iβv$^`4MEo��?�� UOO0t~�I7��nV�%P#�#�"��ܖ���}��⧶2D��K�Ts(��\�I�э$6�l'ɇO�*>�Q;5�أ%�+0.H�p�R�<S�@�󣄕@�� 1n�J��ua���7lA�����B�4^	���<�U��TKt�Y��S�P�.����]�O�V��'!"�����zIq�"��������`hغ�6t+B�N�s�J��%�킧,e2D����c~6{wʉ�+�d�N,��� Fe���h��L,��N_�~��B��p@-yj�+���u���V��z1�fk0�����k��&k����h�N�b���b/m��g�"�jZ)�c#����D�3ۢ'AǓ&���?z���w�PX��sL-f�J�-S��/�|bS�Yw��z���X����w���;��W��u��������,�:=���D��:-��^`*��ֈ-��ހQXD�.4H���cb��Z�U=�r�j������m��9`��|�Q�c[��d�(��������; e���y�Қs[��'��!�ϑz��RI��G@��gT��xpa�E7Q�d.V����ߛ(�ȁ��]���0ߨz�p�`��b*�Ý�M9n� ���V�����+�DL y�pk6u�%?j�Q$�!L�/ߨb��s)�Q� .)?`���wt��.w��ܬ��k��K{����|��֯��M�H��G(�#X�?�<S�9P2�z�ٯ��r�@��s���"�A����
��9E��x�g�������I��8-��L�ٝ햣�F�;��Ď<����f�2$�9>���%��Ch3�f�i����C�)��&D���L���r��TC�0�̬3��g�L�-��Ŀ?'��}�/2�v?�$�]&�õ^c`�������4����۵��Z�)W�e�kꐳ3&�3_���1Vt)�M� 
-�d{j�OΑ�����(*�~4y�e�!B��ߑ�C���ׄ��V�2*5Mྤ=��ĴK�v�V.� ��W�����E�ml� 5����~S���:��XtZ�|�]g����[V�M�f����t�8,��h"����9d�(,Up"#:��%޻[���؝­U����7�1<�*���$ӱ�x������QִWMl�̹�sC(�+��I��"?�����>!+o+�C�mxJ�G"ٌH�PY�HLX��9���p`R��VB������z��e'rB�ɻ�l����{;s�FL;Ӳ�^ACt���I	�A$׮ڔ�uG�Q���3�m��Db����C'�zy�Ewr��N�8mػ�l�x��J	W��Q�p3V���/�C�!sE������٧��P�6"���)͈�Hi`d'���ז�c��U7U$��(�a�W�[�l���/�t�M���.#>�K���˖4e���#0�K<�q?sz6\��3I��%�.1f�Hkt3�>?˼�B��$����r:2���8��bj{�S2����p��7�)>/��7s��Z�&<<�􌄥y�7]��y��Q��QX8X�J7���n6\E�u�y�=����k��B��������܁3/�R�k��!��S�..=�����}��S�DZF��-�F�����ہ��9RIs�2�uY�������߉�0�s\�6�&��p#;4X�����~�/mE���uՙ��"�>��W5m��-_,�4�2�
>�K�E]�)�s�I�8�n<���_ M�^X�eӦ��t{�n0�x?�7�[\��>V&�^]k�������<AP��
����V�u%�U�J�Ϲ�P8�h��G_����+!~O�`{�~Y��`F�6�s�vy���3���5�N�k����	�.Y��L>)�������-!��]�=��L ����%>�F� ]FA(�}h��a7f<��m(��e"9�0ɘZE�%v�9:�v�m�k����F��q��7bw�F�n�M9+�����S�� %���ne;�>E^��k�B?����D���HU�z9�a��-�	z��N]���ɱ�r<�;�F/ԡ��%��_��#�KH���b�r*2�(����e�O0���j+�H����w��Kx���������ךGpJ��Á-��oX['�b:>�֡�h���|&ye�Fib��+5�r�UH�oک�m�����-r9�@��#y���70oP=�wz6J�K�vuA�z�`�O�8���9�2���]�X9-������H����Y@�A�2�gQ��a��U7
��l�q�wWW_��}����Uԇ(����J�)����5|ӇW更�74�0Z�Ǔ���$���� �e�vJ�)kt�ʊ��aM5{D���Zq�j
"�W7n�ڴ �8��NO�nI�@{�R8n?�������,M�7u��эC���7������Q:>���! �x��`���J4;?���S(ѽ�[�~���h0��%�ᯅ)����kx%vN�I�R:�/	0l��WȒI�>,$��������<M���M-�$���.֏��ts�eU'q�䖐�z1(��E¿���&�X��X��w�B���\�����1�5�O�NX삡k��86�դd�y� �����*<��z%P�[��0~vQt\X�v��̔���ҌJԜ��bI��q��6�r�� #��t���������l8=؈�z���]/O�T`�i�,kyn�������{<�
�s�ގXڕ���i����>`������*d|�!K����r蛂�3|��;��/]}p�H"O����kUw�ezW�uMqx��X��ل��
8�j��
����R�)�����Z|��h���	�d��Ⱦ�O�Q���d�2�t8ε��ۦhg%�<��������ڦ꒬����*��ȦS���Ć����|�)�@��"Js}q�C���|4)�8����Ro��ꓐ�5`���B4a��W*�����T^X��QǇ���O�Dp���Ҹy;���s<��6kK��q�!����h_���樞 &Xi	.DOkY��H1����f)KJ}I<�;������=X��am4*Q���&!K�-��t�y���1�jT[�w��,q�)�����J<u�r��J�
�-
ͳ����-̈t֕U�wM� }�Zà�4HnXk�F\Ȑ-�<�i��R�BPxl�ff���ݮgX�Vt([4��o&:_��<U������l���qXNs�q��#+���j 7w�"e]�xQR��'��˞�_�7��֥�W�;���
��Z�I1D�m7�A�7`V?�zpŃ�Lx[bh���w�)LO��r���=(Dr'���E4|�G�vh)�u'1.@��V�H��� U�t�$����5]k�W�g��4�!:��A�0)Vr���8�T�í��	���� �ź�q��4M�>�(Edz�v6�>�F��o~x`��������O��P�}��$�?Ӓ<�Nx��p�J��l��#iአ�`wI�2D,>b��vЅ�)��j��4�h��^��&��hҽ���N`���P׆���ÒЌ���r��bN�*@��0�Z�x�9=X{��S=f��Ż	pŏ���_c�C�p A9<N�s�)�,�)���!g�I���z<
��4E�Vj�Q�f�^}��hC�'9�j�����"�uU���f2s�Y'�ng?]�ђ��Ad���܇�X�b�ȥn���ڰth��߆25��v�>�َ�m�~�d9H,���u���:؇�3pO���g^c�i��X�a=Z5�����s�}�>y1�;�+�))w��Y9��,�1�滄�QA�Qf�P�a�5wt�ӛ�v�R�^�6�� %�i6���F�X���!#��Ϣ��?
)~V�V�����ݒv�L7N(2G�"��_�Z4��˵ba����n�i��A&ByB㔍\��L�]j�y�6�\m�h�V,�ӛM�f%�>�>
2$^��܊*�^	�'�4a3�[�җjFȤeȗ�0�P�zks~�Dr�⵷{v�zא��/�������}H]��;r �s�-(��� �d�hY����ؗ��.)�y��9�J�5���Irg_�w��l]9Ѭ�#!��dT$��n�>��l�xr�7�_�}��V���*����|!nT�$g4�Ȁ���k�6���a#���w0�2;�2
���J�>1��]#&���.ϣ��դ�[�\~��~MP�zt�HJ8�hϋ�FI�����Zy�'6|9xS��^,eϲy*�az%�ұ[_�D���e%[^K��v�e��U�����=ų�˪w�۬�O�2��p�V�9s�Ή�6��n��g���35YI�P����/�j8�u�/�\��]�E�/��ڨ#�nj�z:��ʫR�}}|Ț	nZN��[��(�+�����6��U��
�Cz����t�r�f0g��[���󥯰���nx�#B��ajT1"q����I�_%'���ߖ籈��v�6��3�!�����:>�T��"�E4!�'��Y����T�ޮ8��Ԣ4�# #��0���a���"�7�D�}rBB���Z7v#��)o�FU~�X���k��c��p<��v�@�kޘF�C�b�%�����/�A�;��EK�Y�����~k��װ����2�����r�&1.�2:fg��b�/��ڨ��2����u����ʡ�\&��jj5=2{�g�S�_��6rt��#C�w�ڃD���
���(�P#U%V�
�9��3iX &X>6[��7'נ �{M�������g�F�<oƜ�A�W���}�}u3[$�a�$�nZ7��lqj~ 3�ȶ��b�S�An��e�_3�c�%(�G�g������b�M9C����,N���q��o9G�6�O��a�S���_X_&��R�h=ʣdhg?�,�VҿA/q�����/�� ��0�c��Xz�D=0I�T��8`g*7I���H�_'-�L����Ήm�a]��:y"��>6q��o���n��Yʏ]�'�e�]V���#��/��˚����Vk�A"��zߤ��J��	����(@i��������XaUE �����;#�C��˴��I�t��y�~�߆�7���pA<6c^-Xa������T�o6��eE

�r�7��t1&{Vߗ��^G����z�?�}��r�⅒ 4L���g�[D��iM��tTx �7�f��a��8�-i��-�fǃF։f�<���PE��4A;r��|U��5L$��m���E�	?;D�I.��5��*\����&::�AX����R Ar����[��>=®Ʃ9�AE�����Z��S��1�ť������ W�ǡt�J5[5]���ً��F�!`���y���7�	l����`���k�˨�#/b��[��,��dΉ���&�٤Y;��l0���>�L 4����]�靐�{�l�����BC׎�0�0��]~�'a����\fCcm�Gj���9��K����]-˼���v'�������p�2k ����f�}� A�O1�bHP�K}�cɽ:n*���OJJ�9�v���-�f�6v�!Kg�@� �@��qƨ��q4�sJ�lT�UTq��R�r����:�/����G��TB��f���L*��9G��(*���Ҽ���]�(w��+�Z��gF�p�kC¡�n�ٍF��b�}�-�k&8�kC��!F>�I�;\}��NrOt�Fւ9�l|��e�Q�lo����&�u��i�˙�HHZ�:�Ԛ���#�I�Kf!hѽ
ՐIȹz�<\ث�1��L�r�⦊�x�G)�b�]�n�!F
���ya� �?Ӕ��RW�Yyy�b�|�њ��̜��i���7s��I�m�v�p��R�
�x�4�%A��<�0�x�>>���YX�.$�����'q���wm� U6q>���5��v�~�c)���Q�L4�'�U�>E+�=U� =����$���f�&�l�%�	3�#��#������`���m(���A����;H�RWO��z"������*�E�X��vi��� �Lm$��i�a3s�ڤ�f
01����V���w�����O�4�۪�bw�( �Ӣ��ɞ�]�I�IHn��cr� �e���������׷.-]5'@U��=�l'"�;�
�|M�~ϴ:�ǉsf?��(B�Y�d���^RY0�6��Qi�~l��Y/��Ƥ�bmM1�'N$@��ڄ�2���^4ZO��H�H���%���B/'_&�x�
H�!㿮{��|�J/gn����tW���]�,��W�y1�<-٤B���#O3���Zk�Xז@xSܧT�4o9�3�
�v;##T���"���e�T����b�>jm�N����M)���D�����ӶO��⊒~��A@Kq�dԵ^S��e�thsm}5��\��(.*+5�~�0�f�?�2O8�� �'�H�9�;�)GU��ɴ��(2�aq�m�Cͳ�w,�swnăЁI
���YC�ؖ/
V��Ǩ������
M$���ac�I��4�C[Z}b'�5G[�^�Ƹ.�������8��t~��}L�yڂ�Dt��:
T�(�f�
���8��b�P@2�Q��/C���v��)��
l櫝�����`�>��Y\���Fm���)6,{#־c��/\l�=Y�K��K��_�l���M\���$�n�/~��/o	�d�C�&�$}���wk6�h��h����L]p��Mc������?ij�A�bſ�M#Ti��Py�kJ|ި@��g�vX�#1���J�Z@>S �-C�R��b|M�G������q��1'���	�� �g2DǩK|D}T��/�FCu�h{c"ND{�4?��|j��ziꏄ;92 4��L��L� ��6�2�3��;��no.=K`*1N&��zڨ�3�Жՠx���\g:Ey���	����X�,X�}��Cᡩ?��h����rj/�)���8?����X�}n3�{�����V�pkӦ�o��Q�%Iff1!�Ί��R/h���R��4f�N��a�R��PG 깈x��9?��]�mC�qܿ6%�dK�Y�N��Ts!�a�~���
��V����Wg��R'&\�����b)�s���q0�g��ܑ@�f;�e�$H���U�^���C�A��_��Zr�A���^���̣�#E
 ��<��6��V�HJ:&�OJ�LRG�${���z�fW���z�eq� �e�S����'�,	~�re�ې��	��І����}D���A���0�|4m�� �^%�H�t6��3���(P��Zf�g���Z\���D�kX!8��n���8i�ݓtH;��YW��A�����i#�?$���֋��8���Hk�9>kG&\�����Y��dO��0��(aqR��F�3��ao:�Qzʔ�/en��T��S#���5=�R%\�E�G6�J���q =)������x����=�!�
Ќ�0�[�lUj��x�ok�
��|s�{��|�#H�yY<-�E�Ȍ�n�f��9|���,�_���f����w\C����Y+n��$�;gw-o���R&ç�=f�:��!K�_xҽ\S0?��]�׸-22uו� !.5�o�<\t�|�0��oY\P�_��k����*肘�m�ꆞ���c\�r'm�%�L��~2�G~Y�6�~ƚ���=����	E[��#�9���z��x7�����Y%��6"׍ʛ�2�	����5{3%��?LS䀒��?��Ptѷ��gRT����,���YnZ~Q0%�U�`'NmX_	��f�R4�&�����Y[O�&]�s��K�`e�F���5":��(��;ϖ8��1;)�'�����P���)q�]�l���c�s9��4cf��I8�����
	7&�]�Ϋ<eV	 �./C-�^�9~���ۀ��q��T�Z7 x��8��;A�B�!����+��mf)�zao#���6���UD��0����?��q�@� � |�P���Yb]~H��Z�*?�\�������u�K.;�<#��9��K�� �t����v�:�f��;�'�l��+f�jk�]�e ��G��1w���nh74�Ք�=i�ٸ>q��E[���J��:{ܛ7�Q�0�!�L�*s�.	xM%E�� �c��tC���L�N�v4u帬S�U�7�.r�:d�?d�爏Z���0���i�#�%]��ZG4i�#��,����mja{u�WĻ���ɐ��2X��5v�Z�����HJ���䢞�$�'�@�þ���$�6�4ǂm�������Q�o��΀��t�������ʵ�DɁ` nOrh�Ԝ�C�3v�ؽ���`����j���\�M{R�@y�6��TZf�u�L'�ei�t,5���L�A��Jx�I���O�?��Y����k{5���7��G��@?�H����e���
�s��U�Tg�+#x���CvAݜ�Z?�+�x�n�4�d�8�?���h4���"Z�X��ҫhu}98(PO4pu�j��8]��s[�u�>geP�H��`�v��>��sm���k���S}<Wk�� u�L�I�t9)�~�������T�m��~���g�ܳ�:������˃��azۦ�����*��h��Ij��ێD^u�8Ӱdm�N�Sml�<�K�~�K%�HL��"$��~<Ϧok��j	��ź� a���h�Dry�<��\�U��Gj(����ә.���Sll��+�����`�����kVD6���̟] ,�~���wr�F���g��5`���L�(�������!a��{2�VA�����e�`�����t������}�~�lC8K.��I��,EswSy���Db[B�f�5��u��e��vZC�^o�x�-�� ��-�5:w~i_��E�F7���a�� �]`�W�2b��y��RJ�0���ĕ{�ޔ���P@�CɊ�Xu��<ۍD�*L�q�s��vR?���
kvt`��i��HC�2���䆠�:��N������l�N՞)v �L��&>��zj���Y�Y:[?l_E����}�M��}��0d��"��e�c��T�i�ž����C�"�M��F^t�w岧�|���ߘ��2`ȍ?�(m7 ���K�TA���y�]�b�)2����쑿IQ�����}�P�?=�W_Wp�@v�8(�"!m�9�kc\��K����K�e�
!f���$��"6��ǅ|0
E�ʲՕ���J5V,m�ǽؽ=c������u��/�!s�<4��P��b��k�9�^Tk�l/���\�B�N�,��J��fD���߭
y��u8�K��&<�ǣ�7l�RS,��yh�H�#Ǭ?y�ITݎ�V���Q��@��k������ ���++[�b����'�aO^�
��2oZd���
��p֣�{^]�y��s'�Ȓ7�}��+��`_��N�g ���a	I�8�"1��k�K��S����t��2��?g��z��c�xL�FzwO�薉߶�5ĕw]r��8'�(t��
 ��P��&l�5�ѡ��A9ї�<��`9)q���~x��1֥ ��c�T��/�)�]���oqr��~��Pd�J�l�
��q��=�Bk���OI\d�A���t�gR�R�Zy?�ڍ��j-.�����?Fv1<�([ ����R�0�ި�%j6txsV�9�Q���ڍe��B����#M��}��i����` ���j��������4�2�v�p�u�cv3*�Th��.T�k������}���J��Oܗ��f\Qo\,��
uk�9�u�WG�\��)�n�7�C��<r�K^����!��f�������V���5��O��n��f���
�~�'x�~B"W�V�������T�Rr�q�|fZ��!2o���9_�(1��C�@;��*8&w��L~c�9����^������Ŭ�I����`I�x5��x'�Zo�_��{���L/�\��1\ '�w���=�=��v�$���8T(^A�jy�����s9}�LUA�J�� �[kESF+52cR:Uuym���痏����~��C�L�¶f�F� ���Kw�����9C�V�F0�����K�_A���ZH;�^��_�{�f��ۍz�܃4miWY.�X�5 ����SG���:�=�s�}ǳ~�|���[.N�ܻu0��i��Dj-�4CO/T�����.�Vi,~k]�w���7�8oo)R�2󌣱n��&�-�8������`�7��B��cS��)�����>�"�;��7
e1⬻џT���m���焳����J�5���Y�νj@\���7�
�tay,�z��e����xL֭�2�'�S�������Uo�LG�'D��x����(�\�,1Iq��m��z\:��`�w�����w

����I<S=���� <ޓ�z�L9�U�yI������y���p����354+�G6_���\�s�
5�C �~r���Xu�o� "�t�RJc��rΝ�<%ƪӬ������p%�5�QM�ڕZF����"9~x��m��@�C�]�b�.��
��ʇ&�FH-�F^��r>���]�
��s<bZ��[�|6X��9I��v`�]�-�	��Sy�s�O�>.&�x�M<����*/�:#7��
�`ĝ)���f�A�JQ���K�T��G��<��1�c�&�^�:2�bnGT0~p�u���?��2愋�*z6D�>m���D��҄-���=���m\l0�GBc8'�Pޘ��Ի�����
[���`�*���N�M#6�87%��1��"gl[��J����ͳ#?<�~^1D̜UL%"�ٷg��ӫ}�<}���D���v����p�}s�XG�$���:���Hl��)`B�#DZ�Q׼`�Q��(B;��G$����'
i���U%�5;��^M�	cĜ�@g:��<Y�1��|���!ߧ���$��/~��+����Ӓ�2cHd��;�xx�n��	��b��tT�s�HTض%ī �1j�t���3v�w���1�9�q�����L�4���e@�aXB��FM�&xO�4�>�TC��l��ȴ*�)�mW_������UbZr�>#D�V^*B@;�!�&	u�%J4�,��K<0:�Yj�S܂��r�Ɏ?���}�m� ���V1��Gc�4[O�����T=V�9pz�k�����v0�o�?8�b��� �	*�[+U���5��k�"�]�F�E�4�M|��X�D��w���o4}y�.�������(H��A��;[�X�����SS�n�����1�W�wmaL̬�H�8�E��=�|FF}�j���yiÿ�qv�~�\��#013�<'�y�w�0�v�Y��Q�&�<ݙk�1�r�;�p�g��b�H6�.d���zd�ë(&��K̸�����J��a�Wo�.�~��bݚU��� �<
#�;�	�8z7S.:�y�<�9�����d�\R�J?������woe�荲aV��'3�6�d��x��wи��h;my���;_�}ߟ+�7/p��7	G*�E:!*�Rs��='��m�ܗË�\��n��w��CE��Ħ��nWv"�j�}�NwG�S*;��K���-�V׬���6�7:��&��Km�W^䙁�|W#�v��ۨ�@K�y�~�W/���J;{�˟\#�}$��X�,'c�����
v�A���9R���-�zS�L��GD(P4���eQ��*�LB��w\�ִ�<Z�s0�m�}Ӕ�B�'x��0kW�/����6-�fT�^�{���Q6���DV��Ρ%�B���^J�s�����^p�ft�1) F���o
��a�S��faY5���1+���A�(�4�CM@P���Cȇ�JM$="�ʾtw咩�J-�����(��%�G��2��-����>I�}]�\�py��A�,�a�º�z'�웿�3�=�*�ƎE'}6W��C~�GG��a�6k���\�^|�0w�� �S�$����y都� ?H�f���R��yi�y��r�N�K�Ĳ�g�.����g|��q�_�b��`����d�R���Ru�F?c?�ôp ᒒ�RX����5���_���̑�@f�p)�(]7�S�;��ʠǞg+��^�t���n)Q�h%x\j�h�\0��	��?��M߅�|)����&�n�K�9�$Рz+Z�AkJ�Vj��"E���G��F���]��������9sUߞ3����G��z�'C����A/*o�W5W/s�r����NEYY�җ WG]_ �W���J���*:~�q:�i�u�f��:�>x��$�pR��wh_Q�(����Ggd~k"��x�ϲ�G7Ѕ0�'��QG"@;�m��פ,�Yᳮ �����#H�L��/9�4cA�#�6@f���t:$�Ǝ��R�!��,�>ǚ�X:��w��'�=E�TX�3�׺�����7�.z��%өi�K*'�A�`�&�����3�q\M�b�P?�TV36%T��"��NPFs���N^`儎`���Q0����b� �����ExW�[�n�FBׇ�M	+����e�&�F���a�}04q�x Z�L��w����'��Imo��_[1�zM�bL
�zI����A��$��f�)l3��%����Gw�cR`�_��!05��7�k���mt�����)��w��ڐ��D;���SC�2)5p)�|�TE5CtD�#��3(���^q]���OPL��3�
1�6��)mR����ln���JcS�]iǣ�TJ����T>E��)/F�3���Z�Κ~��s�.iZ>}\�1R^
�c��t���frY)�HF0�i�Sq4\��y4R�N�&��|]U75��"ʍ��Xߒ�
�oIX{�
������\�B�g�&�NXu�ʈ�b���eJo�� ��I:��a�C;���">MP**��-*y����JQ�����S���='Z��TwUα���X&����l"�"w�R�f�guy��?�6�j;��S@�u��b��1��4���\���rG����=l��b�2 ?%h�P�K

��I
��A�`�
��_]@�آ��ÝH� v�M>x�r!*v�
O?��9������v��
��I��������J��V��>~�rh
�o׀>qd�N���a�<�pw�c)�s��I/1�眹~Aҿ��/��h0�+���6��zfGʘ�@�]��g�<ބ�^[e3��#��Sk
�7�c���VGq�L]��&�NuR��6KA���w�6A�kM�����J$L�Q����߇+F*�O+G���������u��!����"k�8�z�C7ְL �~��Eܺ��E�y[B�}�#��s�`�4F[��#����4�t�}����teSy:��= �m��t �Ж�P�8���6ux�Å��F��y��ttc V��a*�2�.8i%:����8��3�!�'0����`͆���V�nQ���W���P/y�yp� �����a��2ߎ޹�C�H�f���h&���s��d>��h��җr.4J"i�ӝ�~���/Z#ܑ�g
=m� ��u�d�%���(�^��k�)��E�VA}��� �N֢BF��#�$S� �V
é�5��G�ߖ��~��\�⁏��߆ڝ~�s��	S�D�����˥�3Y=���Cx�ž\�b�|��"zXz��j&Y|`��ޟt366!u��CbZ̴�d�<A;[�A�>�p�أ����� �f�4������!W�'�#�+&��c��E���1R�a��|���+ڱP7FW�����_u�m�8���3J^7o�5h����St�������\j��v��'�R3�]�������S|X�{��ҙ��ь���Y�����$�j<�V?4�xa�Z{-��B��R��������+�t^��Bc!�P
�z��t�ѽ���u�����D�3!�ҵ�=�&�(�m��MwM�*-9��Ϻ�݉�v;����&6[�m8]r������{Q,0�e9��B_3��'�ӉSSM�gzH:�|�/X�E<|�B\60\'-E�z�yg8�q͂<9	�ZQZ0}o1m}Y�\��v}Zʊ�mFP׳�@
��X�_�A��~�_�w��I�<c�=dy���L��/�R=�t����k�rQ*(B%K��@򗋾���E��3q2����~e`��9��pU��)���~��v�bN��@�d�g-��5L���#(G�9R�s�����LK��Y��4}*��2i��s/��4Q���W����;�0�Ҳ�Jf��<P=ae���	e��<U�ʒ?��@��BP�C�������\�ư��R����H>��2�q���n��o�N#L��wam�C��A�#�C���^7B5��b�J��W�9H'���7W�$)�𡦢� e�q��]AD��K#I�"�	2+������)�������;�L
cmg�)��ҩVֽ	/�Rw�{������fE�3bf���_��@t
��QPj�e�ۥ���fw�d�R��K��8<fF����+HP���շI]���\�%wn!C��T����9k�ӕP�o��,_��1�rW=����i~	V�2�u�Ą�1�B7����ɕX�a��堤n�lc��g��)���2*7yDG/��)�t(t�S��z�	W���l0$���dd�xy,2
�H6ALV��!�f�uS�<S���ќ����i��.����Ĥ����8�01�y�_1�+
Dv�k=��#|@2#���������$&!��'*����v2P�N��'��|��E��v�lJ�מI�g,ă�V�'�BR�k2���*1�=M�b��o���f�	8����,��������89[��_DE���ВR a�0�R���:y�0R�%�Vi���F��ǅM��f��M�������k4������+W-Ї�����8�4�@�\tQr�Y�e�ޱ��	�"U�&��Qؚ��`ym�cE~���-��oB�� A��w20��Rt�d-�7U ���	L�T_��KE;�{��0"3y��z6X1�P�~A9�M����v:�>����q����r4z�L
�#2$���{�D�GS��b</=7w���:�G[��sKH?�SdO�܌�<��IÇɹ�>út�ո���[�!w�`�4��%�����Jp�vS� ��������_o]0����[8�ِ-{���S����N�Kj��Ȗ�Q� m�� �TC1~!B���exǃ=��o��	>�(aW�1J'�OF;Pc���ϔ�φZ~�;.(�8�ž�:X-%��Zm��e��N��ƫ���j K��a;fN��� �b-YDb�6�86�l+�ݫ��y}��g����Q�"D?"���r{@��t�my��f�'�Z�����:�}����K�� $d�beLiǧ���
�
���J�p��6HD�q�l�A/�����A�%��l3j��M�k��W�7?��w��x2�ɯ���A�-D͙����T�u�*�b6d���'�I��b;b�[=�6?��^����k$��{���PF��nmo������Ղ�f\��������M'��������d�<l���,�݉������G�hk!ö����&�s���MF�������C1��N�,h��5���w�}C���G�����r��+\�P�9�n��^�.a��Eԓ��� �x#M�<������h��͠J,yqE�Pb�4M���X��c��)���^�[8Ɩ��~���R�����=\ `�_T���,�m`kIR�Ł���ŵ�ۓ�"S,�@����B5��g|^K	傧Z�*��&���b�ꇹуw�i����x^�F+�S�N��6l��=qJ�;�b�`z���	|�	�v����m��nĒ��֙]�L��ԥP�KRS?�ӣ�m��E�\���8�"� ܿ��(L�[͝��aW2���ٺ,�Z�_½.�:��2~/n���]��٥���lMX��Ʈ ��&�Zϱ���Q��gS:��jJ�������J+9yW����/�l��Ч����?4~Q%���*�$>�Y����I�P���7I���@~z+=*�˃;���9��A�[�X��D�;-��P;Un�8R����i5��V|D����ZeY�|��z��ZsB�/*c�o��:�%���Rg�#޴F�f͟x�����n���E�u?�X�_�E�iJ�~��c�=eZy��{J�m�4 �����ϮU(>�->>���Ɲ-�)k����g��|�+e���טsޔD�̈́�w">��
�M�D/���$H��zj���-���ē��1]��D  �ô�}.��PO��a,���:��Z�f*���l���G�&�1�]Q�6��`_��_�E�D���
�r�ѥ��$9��[�cϤ�Y�)�b�!xwg����?\���U����ߧ)�b�֌V�q�s�n���G������T�s�{�.�L�]�D�s�FΈ��^:�9��ۺ���w�����sj^3�\��[��\�V�������BG0�m)t�K�E���K�Z����(]���fT����1�
��c������������74����j=Q%�k�*#�9�ݶ����q>_����QZ�8�#7�����)rȘi"�!� �	�V���h2���'l�����<m�� 
捞����0Y����)�Z��q�$lQ��gWd����W�QM�xf"�
G�,gP�T�N��I咛��g�lsnOd]K3��7��m¯`���,�m�OW���^C,A�������_'/լ��n2�����g�_eW"(Z(}PE=/�g;"0����~?�L}vy.6�q]r��|���$<2e)\�Zۑ<͡��S��T��S/&ԥD=�;�����IwA2g�P|�u�������%oY�F� �km��!����$A�-����Ǝ�$�sa�~<��\�_�k�>mJO(Hv��V*��#Hӓb���L��'7�aE��rǇ�$Ɩ���m�������s�-@�|h�*�{�v��͊��p��Ƹ4���:MdQ�@/h�!�e���[-F�c<�D�2J$��a&��U��n��r�C��{m���o!X����7�=��Km���\���J^�ȳ�(m�K��S+�?f��`�>FWT�/z@����h��䗵 �'���<76�_3'=D���C\8�-�tsm}#�#֪$��K�鷻��gos��`�֑rɘ��D���B�a�]rej9���	mR�@�/ka�>{uL�eE�����&ڤ��T݁��4�w� ��>l�W�cD�Z��><Ȗ�����1?��:����b߽s�AI<�s����`4���m���%��.�h��<����K��N��T�&��^��+H��|$
yY-HQ��Ϻ�8������@S3�A"vT����
�h�~$�ML�a�`˔@�G򘳏ȟ���w~xuD�Ҕ��t��Mn3e���R���M�(�9��@@��"�%��/��@'^I�TD��D���:j�w�V����hw:���{��^��PgL�1��ʈ�N������&i�Iu���g�(��8����;�l��k�5��֥�*�a�s��)�|�!��`l��e����PB���|7�)�̼c�Rz���~�wF�vƑ�}��OJ��i�=��	a""w42=���i���!?	�wVN�{�;:�"0�V�chwv�\7����~�W�b��=�eͰ�� u�U�P��7�1xV:k��%`��KƳ:$��b9 �?˯��<����&�y��A���TEp��ki}���</�-q+f���O�҃���B���%5� �|MoJْ���X	�e�c|��d�p�����W�c{&�L�'R��r�3��IDa��~�h@r= �J�lD�hҹh�FPu�YWK��e\G�k������×���{,�}յ�x'Lb�����/j7:�_����"���0� b�����Gj�������Բ��D��ISO�OZ�B�Z�][�Q+�+�����D��\=���V�*͔`���q��'=�AFEb��7l�8���L�B�H���,��Q���
�[��HnSa�5��f-�>�xL��5u���RY�.6�s���ۧ��Q$_����a4���,�UD+!�@˃K�������w�\�>���.A(Y�r~u4�f��/� �BU*C�c]���Bt/��!�#�
�a��GϾR�VW�ĥ(�XZQrJ�C%c�ʧ� .fިk�(?^��8{CW؇=.�F��ñ�!�r��L��I\�|��5��+	�2M�AYh���U=�3�,�b���|w.x��,Y5� �s�l��������'�����?��ִ3H������H[A��6/�r�c��ufcКa�
K.Ϥ��z�'�V�&�A����p~>u��2��E�*�� �ϳEv����禥��e��<v�||�l[72#��@������N'���!��>���YX�"�V�媆�l6+oV1�'�z+�6Ov��|�Жю�V���3�c�&�Y�����S9��H���5pz���i���9ӷK1G�{+��	D�;:~k�=�f��Q�5�N�+e�w��5���c.�91�\��(~Ӏg��?�kb��~�Z�v��!�B5�6�C�f^9@"N4R�����N���c���9p�(yޮ�c�ʚĬɳW��-��F x���ms�m_Q^��!G0��,[���*fr���<o���R5���2�y�_��v4S�=�ސ'SSLc�	%G2;�Y���'���6*�<�ќ��?�hԥ=)���7I���,xf'Y�a����j����d�ǋ��"y/���������O�b�W;��a�>��f���rz�e�7�Z�\�'T4�{�qz�;����>T�~a-%K�w
���${�O�}�m��g�u������\+��'�1�ݩ��������r����֛8Ve#�;���8V؏𜭕�h���*����u����='�ĳJ�ꦊ�����ʹ�u��\	G�e@0d�A�-B�uR��$Aɮ��
�\	y�7^3�*Bڲ60�2h��?���4�Jy4���w�$�Y�7c�X�c�Lzvy5d#m�	C�6����Q4
����q����l���)��]x��[�J�R�*��ɳ��?����_>�Y��s{��=���b�M�9�ُ�["�R�'Q�4���#l�xѺ��-I+�C����T����m��}G�䌆N �nRa!�����g/��O���bIS��E�����G��	�o��[�A�y�v�h�b{��#�̭�beS��NE�¢RBl�ش��b�a��n�R���9���k��A����2T	|۝���L�O�g��	�'ُs9�7�vv!(���k��74M��C�9r��N`an�!�J�]|��f��)��l�Mu����#u�B����1����{,D��p�OVG`@2R؏'��9�=sK��|�z��@*�)B�����n�Oˣ��S�?$wL⴩�g�iE=��%��>��΄���O�l���s��Lp|��>o&�f��wv	\������X�O�4��� f�d��X?y(�~����`v��E�x�g�S퓖;�b�n���?���!�sY��)�V�9�r8�x���Ek��:��0�k��K��c�v��ű���>��~�"� ��d��������͘�I�k�M`�R�[W�j-;5�k��������q�A�\�l>�K�	Da�b���\y4A���ݨ�y�w����5�R�O���%�����D�F�c1qYC��<"���6N����Đ�Ld�0�t���:(&��)��n]+���{�9c꓍!|^�rej�+M���UI�)n���È$ �$D-G��&w����R}:��cӌR�k1k���I�Ig�{�Y�$U��-�h|œ��w�Q�c4�����qn�<\R��i�+�,9�.3���6%������.���oCK�'˛z�b4v�">�s�y�S��s'��_g�R��
)�=R�2����v?��\��K�b������^���Kʍ�F��&��PX���A!���''���-ڔ-4�����.�!���J{���P��}�`CEp��
�W[�_4�j0�#ެ��b�Ю�tQ8N�������_UWQKo�)�@E�"H�u�s1�=�٧�L%�;���D?�DR??BA����;����u!���A �ZEH7&���[�{ZS_��`��'Xy4l��尌��U���Y>�onnJ_� ��8�lNS��g�=�5����
D��� ������V��G���!���s{%��D=��
h�:F��N����F.����C{���ۨ�!��ˠd���W>��V+�k�'׌�ׇJI�А$n�v�N������(��!�ER�Y�t��� v�n�[�����x��Q�-&X�&&��d��|E+�@J�UfL�|��JՑ:J-�3�[��_@+=��$�5���v}a�0�SdJ�冇?�@j�G�r��w"ij��xts���m��N��C��(ż[�j]�Aե��u�lƺ�!H���JO��r�
u�Y�r��l�Sg���	��$+ͧ촣`���"����Y�t���m��xPN�>Wi��?��P�3@L� ώk����K7��R��~eGj.<y��eS�:�UW�C����+�j��M�j5D�*s��%�^Uޤ0�i*
�)B��Q���~]*��*>xW��<�G88�ٟN	����:��c�&r�ȑ(��O:��]���5	����<P��?�����v��g�}yɋ(�ekQ�59Y�W[&U�����Rp���K���
Z�$���/����s�bz�sF6���&�O�`���/KUѧ��1�m���Y�7߯�]Q���7�iI)�|G����^��`�x�����YP�9����X�N!�V���y�-~�q�o�˲/ !��юC�W{���ʧ��k?�	D�`�j�Q㟆�n�<9�3�80yK�@�_��x�x���C�ؚL 8� )"�f�}��RL�]~K��ݒ�"��MX'+=�W;Y������&�K�o�l���~�A�$������F|T�A�*I�f�T�!HTa�|�R��ϰ.�L�B*�#�R��v�)��֫pK`�BF�"MZ6D�qwi�P	F������P��{���'Q����vՒ �"4��V�w��M��� ���Zɵ2o��Q����aZ��������X{�=%�b~J��4���>�������tL��3j�q��0Z��b���Zu-t���1��H5��~�W��r%b@/B3Y���7Q��M���l�n� İ���<��2:2����iI}�Q:Id�Q,
h���*0X�8�zoK/�FɝX?Y�_���V�ɴ���8�! �����M}j32͜�.y�:������;┨�]	EV��c� �����"/��2�v"����v�;;�wO�{�L.���;�E����ش߃�W�Q{	A�Sf�"�Z	G���\��_/�z�!�ڲ����\:�#
v^�1�?�́�����
�����������/��a���k�oi?����|ו� ��T1A���$����Ql������i������EF~�K��0�T"�M���y���aJ�0ԟX8;Q=�'�A�3Dd�/�$�����Q�A�d���d����M_�%<��ؖ.s�G
���k���Yu��a�����O?�����Rw��9�
B7�]�@sCY��'�/�c�܁4����$�12��>3 �z�'e�m���G��.mG��Z��M#`���4e�*A(`�p`ކf"T5��'�:�;w�����O��Գ%U>1XJ�G��7OrOۈ�0��n�m��"E|V-�f�kx_p���NdT��x,?��2'2�Yc��������Aˎ�[5H�,##k2���
��ez�F#
�uOv*5�x.'$d����.�]M�9� ���Y])C/�(a�p�L;f�O�l�����@@�ǈ&<p+z^㖢:��I����#Fd�{��@X>I��{΀�f��e3��=zX��5F�z*�5o���y;R�U�Y|�~��w�����:~����Ъ�`���7�Ə��絺FpIA�N[���j���r�ȼ@��ĊEA��vA���a)�`.G�JՆr�*�{5"_��$4
�f�W�?�޵�ۺ�\��s|�4���D �|G������Y����p��ͬ��!�K0k��?��b,U���@^	�]n�������pP3,jxcz#�����B�����f���,���eh���o���~��]E��jҳ�k�Qs�P �?��4�C���|��d�%bs������Ir�{�t�ŅI�%�0�ۦ�QI��'�'�lQE5E�w/�Q��=�"����]=�	 �eW��b*�	����	���~����CX��vԨ���La�`�7{qUe@9(P�D+�S=�'��ʡ��	<f��Q;��B�+��5GG�����,T��6���������Y�{r,��o�Ms%�s(��F��a��TQ�,.�W�?蒂Y?�_�q�g4=�耓戴g8b��� ���*#y^��	��?��ABcA�B;�by�j�c
��, �K]�۬���]P����S��3���O�*#U���〚%>0����B�a��&�9bS��&^�9{��"���) <�c�c�v� L�-��� /,�IuWġ��Hd4�����	�W ���J`l���X�|��
�U�ݦ���t�|���Z�����P����a�]`b�������I�;��©�����=\R^�l�sFn�2���N��s�0'lQ�)56S�T�.x0��nF'�#.�ن^�d���y��K^ö����`�ɫߋ�hL�H^����/����J�R�^]5��tMU�z1��&��E��'���^d���)�]� l���4�B�}іX���h/�����ֈ�
��\���V
ʲM�T�jй��(KX�oԑ����M18��̑�h�"���_y@�"��$��c�_'�D3����NK6I܏Ab�Ѱ�N6�K�z�v-p>��rP���E`�Qf�� �G��'�T�~��.�M�����������2'���=��Գ0��<�� �3\�De
a����t�gQtG;�������M# L�tB[Ĭ�_��]���l��4�a8�|��y'��C��ЎH�>8�l�,�	��*Z��N����A%0�|. ��(�eq�Z�<���b�H�:������nC�oCx*5��D�pZ�e߈�Y*�	|4~���r��a�SIgñ�'��� O!�Izש��i[���:@�fp?�vz-�l����h3T;��xߎpH���qj;�ԡGkߧ���;�{����-1����A�N"�:�ÔA���N3��*Zd0����PS��e�L&�Nl�H�N~�s�6�P``o�?p�^���$ݘ�(Tǰv~an}q۸U��e����� OG|��KNSS��'�QL���̛��:z�KwlN�y0���ߴ�	�4˖)g���&W��×E��ȼUW&8�[���| jN�;�xs�ʪ��U'���F�-�֑ѕ�-*B"��׃��OZ�#.�В	��ɗ0�c;��/��l��@p�#U3�n)��IZ��IM�vO!�(��O�IE���T�y��Y����$����R�=��>�^�]M���.dہ~��-���GDk���YFy�i�6�*�q$^�z/�u����dp<r]i�x�"yء�:��Q�!���x)!3�.�IoF���* �*�#�}EV�,�.4����[�%6��3:pTȶ���XT\S�+&9��J*�_	\P빛;�JeYeAI��D�6Nd��H:z6[8[�t�񮅎l��ρ�r�<L��(�mа��S���P�������i`���hdR���W�!i��I�Љ� 2���P����f熻�!��S�Cy�f	5p�^�IAՉ�9�Y��V��)F���7>��O�$z�'���� ��&��D���AX�t���Vr��D"��d<�.���5g�>A��J��_�]��x�·gXY��Ëg�8�L���;�=�_�c��ry��60KF;n���:=�K6�m� r����9,�'"�:�iGI:жgy�Q������2��F���iVuU�Fr-�X���#̂�mî��p2����GDTߊn���ƫ�
���3�;�[\Js��R �-�o6]s^ai����AI����L�8=�����6"n�/m<�jjB��L��h�?s���i-��A5F�� !�J�u�}TB1�U�[�1�i����mҺ�x�U������]�p�f����v�U�m�_�Ƣ����ʜ��NW�#f��{�^�"a����q7z�S&���å�����C����"JZ�ȅ|M�E�[%���9}�,,h�(m�}gU���l��؍6֘E˥E�>���bK�C��"�M��E1N��q+��`i��60���,�]Ǎ���c%���n\�k��¸�Vl�;ޤx�
�!��	�3��>tHv�I2�O�<�����Z�n�va3_��S�������} H�55a�P���q����/�d 9��Ȓ��W!L���C��T�X�,)`Բ���xX����>0�,�-�Hrs���H�Q��(��
٢���O�b(4GL�q�L�[��)�"�2�Z��9Ȼsއ��^4�9Z#��f�Q��/G��O��=�6����Ch�Hl��6�*��7+s���3 �$[r!���0�6o�s �!�9ѥp0g?�jg*
�?�Ʋ�&0*S��Q�94w�1Xy~�U��lv.p��|Rƞq�!)��9_<���(�imD6]�^HO����q���1W�`�����in.a3o�m���s��_���?:-[�&��jjL�Wr6H�1��i�}V��;���cnW�}ǜ��5O��%�R ��^(��˛����M�k�u�*�\T��{2�v���=�zh+P��4 84�4Qڍ��4�0���A�arV9!�qZ���2�.�ާ��%��.��ք~���$ Ϛ���ӏ^�W i��;.<�0����摑}�6�:��hB��8g���8b![foK�u�� Er�i��ި��v7�+fu�=F���H�B��>��%r�2/�7���>�d�R��� ^{���W+��6�ᩨ�`eB�7��*6�;��8tR�H�+��,����IR��9���)"y/��V�Ύ	��nH���v�!�"�~���f�9�ήPDВr/3��� y]���D_�eB��F��r2���Je�ñ;OHG�ÛwA��	$��n%�)��Q��Pw�d�?n��Z��w�6=�����S]�)lv;�C��R��a�t�F�J�jx�1�zE0�h�{V���z"S�L%�ގƞ�O���S�QR��@y�,!>��ȶ��A�>E�~�{���.���B��k�,9;��(X�9�_��#��Q�o� �ޕ����P�5$���/��q���J�i6c�l��ܜ�i���2O��@K��F�{j"95�i<&��SXaR?�R�E�Ο�������0V=�̦b�:~W=��G
��	a�b���b:VX%\��+E��Nx�7l@d��N9l�]D\.:��y��dX7p<(�)��?���rb3����xg2�����&lA����L��e��;�>a�>p㮖�Ť%��G�:��Z��,�A�c[��5�c�
��y6&&]~�_��/# ���̊⽡��ye�'
	��,��f5�6��vz��t�����t$�\t�i�C����QD~D텠��F�5x�jek{Q�ծn�1o$
h���Vx�/�t�'#�^A{������h��^�w�,S�J��C}���@s�?d��1`{=�i��E�b{@�1�͜��и�ܮ��abN$�ǳѶ֩$(�:�m3���U�  E�^�|Q��'O�z�ەr��܄��bh���5��΁��[�D��ϵ����
h���;�H0�-JLãBQ\r�^1��h�J�\7�`?]�ㅜE�� ����S���91���fV��Z�9 R�;�h��t��<�uz���Hqr����iQ��q��?q?�Ơ(���e1�h4K���69"_)�$�ڽ�k�ӿ혜PK�bqf�mߤL�`�d_��R��:��
�&s`_?�L��^��I�k��<�$�z&C��-VW�Hט~$&Uҡ�X{ �6����F�"␆j��O�1���U@T���`p#]1� pm��*�<���+U�j(ǡR���Ara��c��O�-�7��)@ ��N~�h2���0����ǧMOy{ʀ~��L�W �� �8a.�ܗ����H��0/I�3M��l�?+���t�Y�i��T�Ҭ����(Sb�k�w�WS��Q��as�|3t��&��ƞѼ�(3��T���ݬ��1���$J�o:����h*���Ш�2��YwrvD`�aD����5\yx�E�&TH���!E+/$��"˶'[}�窘zm�턋Y�p��c�/M�R� f�WV�� ��CMV��B����
)n>�]kU<�!�!T+�(u�����m�Ce���uAl�X�u����*�mb+������k�'N�?���/��_�Rg��kyde}��+�4�$�7C �E��hy�7�����Qz�RHB�L�L�!=�
�BUW��!e��/M�Q@�x\�H$C���B�_c�o��<��gr'�[-{@�_�ʒo���}�=�.�4�$��ʀr�!Y`�{�P�j�Ǐ��W�{ԝ�H߇6{�RcA�g`71
w���-%��n�:��n��qc���5<�X���}�y%_�׸�w+�o�A�1���G)�G�׃Z�ht����JI=��ig�>idio���w�^�df��,BK��X����,\\�(8�ob&S'5��D�*�OC���W���m� �IA�ЃI@Aa�1�iMǘ�.t���!�dpL����-;9����������������h����t�I6��WGg���e�Cm3�֕� �e�7�'�%:=�-o}�iK�N �}����nN1�����Mk�[A�3����pխ�:�QڊG�#�):���G�_�N��]ޯ�x�={��7:{~�������(��� �~Xa6(e(����xV�:�M&�_��MTJ��ݳ=F���=;�@�3p�5�ܯ�]ө��e�.@��(?ѱbq�)�����_Q*����������3=[[$.�����T�|qFf_��W�V��߾�P��Z�;Ыi�n ���q����?����Z����o�[�x
�kP���f��n���?Pos���J����3<8{�a��ޱ���\�a�/�A`)0��h�?�1�Wc�Y"��R�
����J ~�&��D�0�����,C��	�3d$wE�(Pc0݃$��U��r�sB�¿�!|�0�Y3_�J�2�u���V���D )�ߚ6RD��iı��ؐ�L*\U�kB*bܢy"X#^����&��|�t7�4���a�3,��&0�v��#	�(�s[�ܝ��z����$@er^�r ̛���C�a��5CE��Qg�X �^�P':��I��<����;R��~^��s� �V�r�<;���<��)JjSرr�^�Th�6/��a�LFx���wb�s���
��׍S�&PӀq��勺&Y+��gL��ן��@p�!˻��Yq�8��ûi�(���(h�~��Tf-�^8�%!��_e=`@8p�2�B��,�+۪<Zoǃ�=�dBc�Q��rK��\��e��u���?�13d�L$6��4B��6����nx�*� �zY�H{�_�4�I�:���I�1p����j�PKP��e��_s�u����#�"k0�M�R�T��j�wU���@�F�?*�.���x�|�F�� "U'���V��!��][��M��`��v�e�["nnS�x�K�����U������OD��#�2G��hn�B����e[EJ���gWOx�m�%~�Zw��l/*C{��N�Wa����Q��7���"�$p8��8^�U�-��rkV���P%�P�JX&��~�fERe�#��:�ɼʚN���,�?��3��oUJ/�r]x�̽���%�����<q泽IFa���(�⛃�$��hE�#�LaxoW�ϕ�б�`ܡ^�ur�}v����覩����g�����ƥ
޶|��ob���'5������LX�n���N�/���<�н��ិ���=�������i����N�!P�Aͦ�k:��f�(F���U��H<#x3��{��d'W���m8C�RY�_�'��~v�#M�{h���]{�]������ϙ�����������s޴��F蘘n�������@S����xrr%�@M��r'';�QCsd}J�w$/��'ʥ�+1#] ɤ�$#��~�fL�ҹo��> �N�8��c�c�@�7�q�T���ܐ�k����.���a���9�|�`F5p���"��R��к{N���7%�VND�K�!�9�-�������K[�_���*����{�v��y���s�(�S�8598�$VC3%��J㴀@!9��<�׏;�$&�G�t�~C�x5�;����A���<&22Ϩ>�d�?nދ��OK�ݳ�2\�"'�I���q���_�L���' =p�$�F���	���҄���󰬍�f
��3b�3���N���D��H�oj����s|���x,���{�8��|��u-�\�#�4L��OM�ɶ�b���[GO`��Vь,t!�c���bO�2����gnG�����j� �M�\�l�����$�>�v/�R%���@�p���7,�����`�G��}=LHaP�?&j-8Smwb�y"�O�nZ��a�0�2���n\���bϯ�-�.8��<��3�0�y�b���4�T%~�=z�i�w� ������l��I3�U��DB�$����Q�G���ΘF ��ؽ�b�wB�@`c��	�d� I��#kjY_���@x�z�{ㆭ����<��b�����k̖'���$C���L&�X�yZa�?����.��"���;�SR;r���0Ϯ�:��I����6���,�h���n��alo�D��,�{�d�br���/�ގ��ى ��~%�7�W
ҿU��=a�L+�T�t�!��U���1��-ŏ�iU'p�1�v`,���\�F\R47(�� ���>�q���=H�N
V/�l[oӼ��)^�D\ᣛ�$�wm�׻9����ڻ���u~+�����?���6���_�p��[��5UɎ_p�]�R������@Sθm����.�rN����{Z�v�q�O0/� ���R��dY�V�PЮ'o�6ho+�6�	;Rx��ƴ�o:,k9e[��c�����m�U�S
��U��Ę΄0�쥚fƧ���1Fj٢*�u�g���V묺-��!�8_�a@6E�IpҬ�2�Jԧ�	v�S�+�He��Y�	
c�%���S�8Qܨ��e
�|����2�V��Է�����]���5~�8Ep�߮tS�.��1���7g�����R&�|�o���SK�6�'Q_,l�����7"Z<�(������炯vS[��V��2y(1��xO�y���?2�p""�|��3��te��̙����'�T��=��]�Mԫ�4�p�Fd�8�.�zCZO/�t����tIc'XE5'��E���"�`Ə�B
�Ij1F0�o��J�d[>��#xI�
�FRi�P��+I�j��@B��p鄊n�N/�m��ka�3�.I��?���	��]ԑmlf`y�ꇻ��CNJ�"��/c.0�<��N���̶�5�0��Oٶo�b>طq��/��t�Ea�N�G/{y��?V�99�>x��{����꿞b͡�{Й5���Չ����L8��@
I�}�ν�+h*2I����61[c��K(�4�r��k
$Ԁ_�Y��,Ĵ����>�D��/�%�Q����YE�׳���
tO�������]������q͝��ʖ���b�e�3���W|gk�#1��RM���bN>3C���Mn�D����X]�L��#x��X��Ȗ���R>��@ ��v�����㢤����߈Mb7���Z�)��pퟝ��B�<�O�Z,)�AC���vu��*xΔqF.陦Y����I~ǻ�ђ��BKV]0kp "*ka����,�E�1<�s�/��X����/�w��O���ˢYX�Jt$�܇��t�C��h	Ύ�q37-#�z���D���
c�0tu��d�1(@8��~!h#���_�l C_�������0�M�ɷ�=1��Tc��:�estg�ǘ$������T��:�N����k���s��,����_߁��g�Å�_��T��
r�
��z��Wݕb�HU��l��^�j��D3!��b��n����E�O9)ʎ�$D��ߖ����z
�j	��n��`5Ց�~9Ҝi�e�(��fjL����?~ 8�m�v<���^\�m���KA��շ��m&a����I�Bhe����9h׿f��(䘱-��y�"�)�y�r�)�x�J�R[�5zU������{n�]���F,�3�%���(������zn흄�i6ͳ@)=�Q_;8t��1P�O=[c�PR|XxV�ŧ��0���M����39�k�(�=$�1��Rڧ�`,�f�$u�S$"�j�Ix�Bb�𬘒�<jP���+u�N��|w�{����b�ԳG%���1vGNS�4�w?'(�c�A~�B����!p|G�(d���N�NB)�%+�Y��1u'�v��@`N�Խޥ6�'>���Jw�dbE�P��^���%W�hyb�^�<%�ow�"g	���,Z���n�����#y��5���$|df[ܣ�e>[�L�mg�힅h�4��c;�ӂ��=�xxH&u0{ч }�x�����pS��b�?:��3N��5mJc�����Y�7����hm]�K<�9�O	�:z�ǳ����xæ2��RHZ.�U���<����[]4�0d�C����O�F}�U��i˃������LlVD֏�������;�|�3#�@��(���&�4=���zxd� >�L��~�rgs�`N�$<6�}�&MŌ�=2XX���f:z�Sy�v���cY�\��6M2�����j1�GГ�ݧ�"����m�����W���&_�<У�Q�����?�DI)2��"N1��7�a��r7����3"�=8O����8Z6d�V�*��s�{����
d�{[T�̞O�̩	�ٮ��`yP5��H"�C����^�;[�d�g-ppK�jyãrW�w�
�ZG��",������
��h)�m�	(�i�qQn�H��dE���kp���B�0�߱�1������V���m� ��An�Q��� (����L��0Sc��;f��B[k�����U%�p5��)�����U�Bn&�T5�֏��5�>-��4�/�T��q�꣮���!?
���j�I�����{�C ~��ᵓC��K�9�T�ɜ4�h�D?>��8;Z��˞���N���t|K�����f��ݧN��x�k�e��Q)�̹�z�������Nһ2�Tf�<WT���f�_�<.�Zςow�/4�n�&���|��cC6ůaߘf.��4�9�%�VD����l���!����$�锇ЪE���{.�ⳙ���\/1�P��"d���H$��b^�K�[��G���w�><a���i"�ـ� �X�宋6Q:��fn=E�ϒ6���:�N�'<f�X{��xj�y����8���.��$G-a�F:鉸L%h���Z�=wH��-�Ȯ���@��d啨#��
(�3��۝��d�O�Q�*�Oa�O�B3��DKJ�_7�AK��d
{�1<�q��ْ��Р�H�ܒO/	v�e�~����(#p
}Z��Jd�/�f�}���#t,�c���?$}zC�QS� �[j�f� �/��X����Tfս�l�`�y��
��^Z�u,"�����):+������#Pi�K��<kI3�̅��N&���R���.�����,���ݠ�;�QY��c���x;�ȗ��P1���2e��;�t#�����<�W0,��4��
���E���8h���0}�� &���� g6����M�+�I��Psmw{J�s1f�H�'o�D����T�Ih[�d��bXU9�t�WK#0���zL�xS�Z�M����.�9�h�V/\�;%fV�ȿŮ��,�+x¬��Ͽ�0{�@0&�8�#��%i���O(2@�>%$�؋�qs�ǐH��i��6�-\�e:p̻;�AH�X����4<�&�b���'9z�+T�n�����s�;U�@?��3�b���X$��6�Zn2'��v����:g"]��l䄏/�?�*پ;/��l!c�@��Ee��&�D*{�L���A;N��]e*)�m���R�O�R�镭��TJ��&�b�gK�/�kt��4�0e�N�["δ6�W@��d>~'g��4�n���(-�L�Y��00B��V:jU��V��1~&⬘��L�Ź���tt�"�9_�f�_�}��^��!�o�w�	�Z�9S�,�����E3@�m�V�u��e�ǆ�� ZV�4�%?іP1L^:��h[� .$qk�N�۰�?�7`�n��I7����FǗ�/�-��׶�hc)N'ͮ�j��}����e�� a���8b����Wb��ix��r����Q�%��&k����=� C�jn�E��S�r��[���(n��k�G�񭁲p�d�V	6)�����;����JGY_�*���	niB��k�L����/DmqE�扣�N4����!܊DHY���l�Ϡx�	�?�u��ye�;�0T8��7����*�D��'4~�!J�&�^d2����
�UhJ�g�h�h��~-|��,3^/�|L��*��K�E3���8��hq��&��K�����ǡ����t,H����Z�72	={�<��������MzĞ�q��:<���So�\J�3�&��<B��_@Ќp5�V���L�۩G1m�9`�Q[&�����ݓ�@?�k�,O�~�)=K,���w�����uɳv�GW����\=��>=-	<����KnB��nO��'�.�rΗ��AVU����L���}�h��v��:���^x�y$�*��ll� �$Q���HW֖�o��^5?Ǚ�X�3��Eͱ�v�����i���i�+M���fv��{\C�J	fP�����f�MUEO���/b&�Q����8l�Z�{�|�4I������2���u��/qW@��h&֏��e�Y)[�͑�1����j$h%�
-��/dy�����=���e߈�����ulp\R���a`,f;'���8�1��f��lRK��N�GRJ�^��)L� �@�7C�#>'�� V�ͫ4�l�,%N��S���mO��(�Оx�X(8�U��
�S.v����[:C~�>�P;ʺ���2���jQ���a�'�	������y����v]�X�)�rC��v��@�l~/�����!m��T�R^э��j�8�e�&��z\��^��g}���"a�ղq���[�sS���l%c�xL��#k���!��^���"�|�M&�_&낑�@���D�Ѧ/����_N��fZ{t>�z�e�W'��8������h�0 V>T�g���G�f4sQ��F���Ĩ�����IF鳵G�׽Cw�J�U�\؈��A/���E%��ۻ�ٛ�P����nx�	�L�ۻ�Rb�yZsҴG:3���@��h�N��n^#L���\�BY�8Z��y�ȴ�	^�IY�^����X����i:���	�A�=v��'kz�X�V�UU�lg?�'�7`��x~!~�G2hk%��H��/b2�^�R��R�b4D�%Mz�]`ū3�ؔ����#�)�� XS��8�ͩ��_�5PL4��q+��h��
�e::Ģ1\��p��j����NA�5�q�$0�	z��u�r��@�r����,i�䭗��d��%%�F'}�giE�\#���y0��]j!j���j�&f0� ��yv,6�&^Tg��4��k@oa���v�	jj����#{cgE����G�\�/9T<	����{}F:T�d�*�����LC��t��ת`�]nf�*�,��S=�[s굧c�M)T���Ar@��G�����L��QCq�@	�rM퓰_����r8���N������a+�?��sJ���4�Jh��l��Xv	u�=��_�tgL�e/Y"����K)v���/�G�����͵1�GjP��7+<^��w�Ǟ[���D�Đ��h�Y�R�:�Yc�1�R�ۂ� hC��f���t�)��q,@�}��%�����r�tԠ�!+_;L��h_Z3�1��bP]�º� p
E���K�ʺ�^X���a�@�<t�>CC1�@7#�5�2
x���mu�KB�ՁP�� ���� =�%����aE� ������L���@\u���2י����V��!�)w���f���J73��R%00W�Hy<kB
�wcjZf�r˸`^�M�jw&&�NGޜ�&w�<����%�Q��M�ꎛ���%h�Hh�\�;�>a:������-��so�1I��S�45������O�n��E���f��w`)<�{�$b3g�{�HA9z����-�£d8��;GHVr�N�łc�����.�}@�9?V�i�Y^c��,��L�E��?���Ug��5����T#@�i�욍BĶ�8�C'���H�SId���6��q��i�J�I�����w�D�B�%�x���n��*�BR��M�+F��l���<qf��2D����sI��,���5�͟$��8L�z�������� �8�w�6 �?�R��M��O�D���e
����͜�4��<�ઋ7t6�H)�Z�8#��]FOA��Uᔞ�l��+&U%	vr����`����A�tT������s{����;>�y+�
�P(y%	(
{���lt���R-�"�f0Uޥ����.���h}�\U�+=i)`��.�\�\%����֦hV+J���,]���n��,�I�b�cߑȩv�0�̓�f8y�81>�����>��R�4(��S���-��^�șԴaʟ>�k�Cw1Ȁ��W.tk��Y�o��s�؄"��m?�*(��! ���y;u�������[�	�&�]���5�:��󷪅��� ��wR��8"փ��� i���t��"BM��?Ä�O�1��r���l-S�F۟e��� �i{�Aλ�)!-�/HSfC��ꋮ��_F�3�p�����(��5�TW�{�Wk��凐�z��f�%�"xJ'�z^�'d�����,��z��z�r�VaM.�A�Sr������1h��ő��Y#P�Pr5YPf��P��_`[��l�ˠ���
���T��F�F=������e
ppq~8ח�>p�K�a�c5���8�X Gu�U�4�2���r�}����&���a[)G�Ϣ'�`<�}hİ�*"�|�'�)mB����<*�h���R!%�d.�a5�밮�p+���nmݮY�J�A�1O����Q��P�(�I��8�\ R'���.�K�Ī���}��Ҳ������g�G� H�n���Rf�ҹ��N�O?�W�2��i��B y�h)c�F3G�S�7�rw=Ol�΁�(�8��^�ʂ"�b3�k�z��)'q����;
ɮ��҈K��2GP�_��j�#�?!��!����q������Clc���*���1���/��y>�{%���_jߟ���,�;�X����l���m���S~D�}6���D��3g�����N,�R����#Q(�m��ﬢ݋��j�y<��듨����]2,O=���is+���o���U���0�d�<2����t�D��t�ﲏ>#_�Ӥ�r��wB?���iO^;����)A�Z�vh���(�IC��3D	:��Y�8�6T�W�#���SZ�Y/mwx�����Ĺ����A,.�Ǎ��/
�n�Cg�(v��_�=�L�T���5U��j�;�7$'+��H���9��C�<�[����-QbrWh��@cǱ�D�-\�`?Η�[Sk�]�M(�F]��?����D���EHT}���ZM�m@	�i�)1���W'�6�0v�f��� ^(|�G����0xMp*�U���va�Z\�oM����W&Z��ռ����w��E\{�{�-�m�;gi�`��Bo��������:*�B�.�"kn�0���n��Y|�Q���6��K<��7����	Lr�|$�֒k�G��}��Mug�
��IGOc�0�8m/�=���6�mg�� �T*V��Jf�� D��)a�{&!����	��ʔ���Ԝ��?V�OM�=Y����g���D(�h�1�.���0�O-3 ΰ�TS����V�@�I���E�^;�wJ���Z&*��Y�*�+JG,��\@��8L;r�.W0\����� ��߭F�����W�� �"?\~*Q����mÁ2-����s���n�u��Ș��}0���o0۸�~�H�#�3�Jvmj&�y��pB�m��|0nF��%0��dہ7���S� ��WW~��`�����pct֑>>�|��8W� }[����Z�x~a���g�y̵ʅ͌�q�&�j���9�GX"������G3��^�z���%d�b�ĕ06��֮�c=���3L�,������31������卵�MF�`/@��X��G��Q80�9Rz�T�Mm8����p�%��BQ��/���Ԡ�d��������WȰ�L����1Hn�B|Y��`Fʠ8����
�i��@�T�v�eA���U���X00�Y������G�D�?{#��m���	-_��d��6 jsa_�n��!%Y��7B�r�Q���N�,^�����י�Ǳ��f�蝭?5ԅ�?�#}k�������Q�F�����οw4\A��Z�}���qc��]��c��%2P�y�`�!�C�����|8Gx���Y��LD�O��$���u
0��$�O6#.�
z��ӱ粑`4T�JCD�pc�� ��4��I��~�ˣ�!�٪�Ղ�u�gf���Ha�ld 騀�>xNt�����Yn��Ǝ#������{Fy�Ԫ�s����Y��`��_��[�5^����"O)��QBe�5-Q܃�O*miS�b���*mI~���9�O��9�l#UV�����EŪclU���}jIa�O�� !�Z�Dvm��D�egEj����D e�.�Ü�iw�-�*�/�c�����w�Ҿ�1^�z|�� ���Ӄ1�ː��X!����ض�z}��>��][/ע�-8�7���6�ǉ$���<cMFtQ7���`�?��k�_�I/��y�
TW���{������.��=���8�a�� [!4a�NP!��xU�#�:ı�L�`��ɳ�I����'�NR^���E�!Y����{�a�Ϊ��}?��	uUt�"�9[��l�ݍ^/���Gu��A���`�{m�oH�� �<�/���TZ��Q�j���R���XB|�� ݙ�A�z2���}�(�a�����>�'�"��^�*���c�I��?ns�m�Ԝ�=N��e�(k-&�Wd{=�[��"͐�p"�v}��%��E�'3� �Ϳ����eU��B�=��O�֑d:FzY����bw��&�(N�)��^k�+�KF����SC|�������)�݊���*����P�h����2T2�������'�O���ƙ���_����<*�9^��Ą )���u���Z��R[G��С�sKnSxRc�~�8n��$e��ߥU�Ҋ���՞��ԯ�5�l�@�b�i��GB5�GC��:���>�؈"��<����ey��M΀p
��,�s+�܆��,~�ˈmuà&DC�H" f@G��J��\���3���� O��Ν�r���ƤV	'*9�Ä~����揆�3�$1�.��R�7݊}�PI|���T����� �gȵ���)|��C���G>ۛ�yI��6�O��Dִ�X�Cd��FBo �i�Գ�I݆)�g�@	z�1oZ����1Q��6j����%�_R�^
�l4��*J�ɹ�������A~�d`��B�~1��ͮa�&�Kg�������M4��������(?�f�發��M��"��~��c��e�^_@u�^c\������'#��.uX�E"A0	w?�e�����SW��Q��M�O����	/���J�5k�����0G�J��nXfW'�g��R�wu�*/��ۤ�p����6�+� dٹ���/<z#��?�?X�u�`��)�<��`�%rI#aM�=�@II���my�a�p�nxp!9����H��Ψ�u�È˺�t�W�CÖ6pI�y��[�%%i�Qȉ��zKT��;�>�����C����0�~D5e�GqK��i{���/L��> ��H��p�\�C����B}5.6�Ҳ�B6V�*���1�� �a6���zN�!�"�c���ct7}Eʙ���U|K0xL�w��O��p^w��l��^�\�fe^C�	��"���D����+5�
�,���X��V�Ͳp���L�J#Uv.:�?ЅI;P��_Q��̚S;d�Q�>2�'��ypZ 6�޼S��
t��m�Ƭ.�f��ۺ׆�i�