��/  S����3�c�ub��_NЀP���t�,ï�!U;�P{�g��Oj*�x �*�'|�N�Q]/];�h-��T���g���X����R�X^U�~U�x&^��֐���>�R>��uF�c<�cp�(�H!��7,��,C�:�E�{G�@g;B6�(��Ov8PG�<ÚQ�9ΚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0����Qe��-I3E����(�l�����<r��R7���aF�:�y��{�v�L��$�0������l���;/��e�|^��<<B?���D'�HM
�����a��R�d���`u0���C��V�4ް��ę3��dV�'#�`[�n1�|��HC`����,���B~sO��5��!?�Q��^�#	(H�?x;��>��^��a�PD�~{�F\`�V�b�:�Z�@J�q���$K���UÁ�K
�y �Y�90y�ˇB�V:�P%x?�� +'�ćx�
�d�(�`C� ��C���Pcmq���jLJ�W�ALOIc��,K9k�� �(7������3<���"�'����?h��OahAu�i�MXYm9���W�gA�"_��XxqY��JkG��R� �sw؁�A���5����Z��^s�2<���̏��Y-%�/���޻�s�06�_�V��siD��x�
��h�t��u��:�b�%U{���oU6� /�8x���d��s�i��x��������)�D3{�i3��*m������y#�G��}�UI�*}GI�P-T�SDP�|�t*}1Z�h��Y��U���`)u\�*��
�V��m�[���g[/�x^�(�c���(@�<Htq$�9�� ����cVw��}��yz���%�٤o�����f)f�$6`��@A����t�SnP�h�7���� �k�N*��c��::�=�8�R��V$�)�U`������t,M�	������#�_m(+Ы��PO�@�y�eN�b�&4�tc�$�&�1���ƍ��B���JB{X�Q���i��ߚ3�Y�@q�$��F��0�k��{�#���q-�	��u�G�s�9>[1�H{K����|Xޔ����ϭ��课���&�jSP��3E0g�a��T�^Im���L�uD�,��.dڅ5����!)�*z���[{f0�g�1+n����H���D�%��p����zD�o���$N�[{(�wi��:�ذ1���Y��i�ѐ^�+ґ���uwy`��]�,y2)tH9߀����V[�&�,�Յ��t効'��2�����+/C���:�?Xf0�C�I���MAĸ��F1GG�杼]VȽ9���u3ud����U2��׀N{�3�j�L�Β��-���i2΋�W��P�GI�H(�l��Bgj,��4;�t
K�aㆦ	e�]���M/���^:��&$��x脀�*���r��)bȋ��k��� �#��=L�-���I7o�#�i첷�{�"�Z�_����ta���J���@SL]�t��~�t����Kݑ5�J����}߂ٓ}r-�3̮�n�뭬V������d������]���������']�d��X:�\If�'���{s��xJ�~u�滽���k�{5,�49�M��Sm*eeD�3�S�Vb_�ł��Ytu��v��)c�i��o���wh���+d�����y�?T��2D@�^*Z��Z.���f�
l��P� ��͸4n�L�Q�:Ciצ�E�M��<7o(j��e�����)lc��{��7D"|��jT�o�j�����\a[N���f�5ۮt����E��|��~,��3W��:�����2�V��~�<yK��������L:D��;[vP s�@�"$���Z��<�v��l��&%��}�'�"�$O���_���z=5������?.��_Z�u-Mf"�*�=!��J�Co��k߱e�{�`�����]H����{
���L9�H�x�$v�!>��n�i�O8lI�X��p"Q�@$�p�A����|�gk�[#�0qz��F�*(�$Ft&���D J�����y��6�<d�tX�T,�^`�� �s��vCOTaRp��8q5����@&p"s��̦<�T`0�We�<֍�X�������6�?����!�����+Y{��dR���Hx|&��Cgڸؖd�m�n�к����ep�g�I���j8�[���j2�x_�$��f������O�������Z	� �7zR�hݠ���̓�h�jX���gu�s�7/e����~�h
�������D�|S]�J���Ñ�x�bW*�(ߏ������}��S,ݖ<��{G��y���~��7�NW1��5Q8���˘.���'f5��oOW�0	�M�*]�T T�ɦ�bMT�-��q�ne����PQ���j5�s��V�>���0��-�w7��3���
�l[U��Իz�V�n���#JXe���l��BRW�tH���đ�z������nq���?(T���o��p�0÷e�&=�&����\P��Q���l�daM�:8��^?��1;�qc��9��0�W���hrzQ=��v�����"�{(�����4O����ּ
��b?�+]*���F�Q؛�gQ��[�e�;H~�kOb� ��Ix�/��k��񦩅,�=o��@��7�*���QET���<V�P|�@�T4s�-�C�?���A\�Ѿ�`�]���\[�^s���:�V;y��q�M왚es��t�Z��̯��ؒ)�}I?ٿ7�@R,r�+?��9�� qEhEWqm�����r!v��-�#�Y�������<�~5#Zn��A�"�Y�e����֘RLTс��y�|�S�'�a�I�px��)����e˓��H{y�Ŷ�
9�8�YVz5��6F���z�f���A��D%<3��z�.�(�0LO}3[�k������P&Xs�_�k�b��$!���7�ƫ�]�nG7>��j1٦wπj���q�"�A�ʬ�_��c���PjK4ݛ�����H(������OS��T�Dohc���oR8���ÿ�X�ՖH�6�#��R!�[����7	���-�5�Z#�՛K�i��#&R��y�L�d��|a�1���|�V.�w�-��x��F
�]�9�ȤW�uG5��Mf����$m��T�jy�g��BzY9-����g~��!������7�w��"�mIX���m��halI��>瘔�>�h�X�kƷ�xT����o<@�`3K����jE/������et,��`�����q��v�D�Ⱦ�@�8;dc���K���N�#�U��[.y��<hv��h8D<����r�,u��A������fNN��wW��!��ۉA� �K��	ZB;H)���ց������}�����̼��C�� �ƻ�K�	�*�0��)q�N�n@��V�]��B��SKJ2 Z~�͘�/9���)�6JX�y�����"M���$��sD��it�ВM�� h������`��ms�]oT��n;�BL�%5�N�7��Ew����4��$C��;գ �`3[��Z �-�d��d#��H�m���ZDbT�[IoPs���]��K|�HA�j
~< ��Y{Z���d��%�{�Y�x�9$�)�Ǣ���NٯS�+�4��=gp������Ȗ�W"�׽TD&=c��,`��f�Y��'S���6m���;�/�AX{-�i��t+��̙$�" ��ʬ�h�Q��aȠ��[g6�h��n�]U��fR�rK�п''���'�4��9��f q��t���5�\�&a#��&��cgm=&i���h�-�u��u�����p�P�b��/������v&\�g3�3~���WP����~������E���-��x=�D�O^��iel�4�]s��uz�Y�,�J�g�S��m#S�ޟ��΂�?E�D&{WAj\°�o�i�*���\Z��s�G�e���l�1ǃ}���Q`�ţ3a?��x�,�{-c��eO�~
�{��N�ĥ��\�I,yaQ�M'aE��d��ߗ���lytN��1�A���`2��Կ >���r1��z�p��'A3M��B
t^��A��~���#�*n3��.e=�:����tY�켹��iC70�?q;n;e�X�º(�����,�)r�Qs�XB��{�c��O�afpx�/-]A'�bX�|eKy�Ԇ����M�Sb�M��,��}]e��.�0���EP�x��oHFsd�z��+�b/�ҷڪ"�[r�:��f�Z�v&����%Τ[�m�����ӛ6`��.���w!6X�]T֟�y����Z�Y�ka�g!�s��$�h$�^���63���b@��	��jk����be����"7 M���¾s��g���i�}/����NO=������	��Ϙ���ۊ	���?@Q��#�t9W�-��h5���!v���n�0�̲y���O�e;l���i�_q &��c۞�x�U�*��S����T]�r�B
�-�?������J���N�|� 5��LK+�y��,?�w�7(ES,��J<�1�Cy�{��3ٳ�:*�N��ѵ�dJ#���##  آ��l)��[:Q�'�`�_�Xa��-R�1�LX����KGs���7Ѵ�$GU�u"7��u�v���:�s�K���SM^�Tm{;�[��E��g��f�6��}cud��ۡV#���<�ָi�M��Q	h%��t��<�:p��.����_oR���~���Ѱ�/�T���L�ER�/:�f�A,�8�F*٦�Uޖ��i7 0g���#
}p^A�σX�ԝ����\&�����4W�9�X�&�+A��WK ������?����}�����մ��  ����c����Ma��Ԕ�1V�r4g9nѯ�)�g%ߐ��u�ey�b�ñ�}���J�⠟���C�7N��la�\l	O״5"��EtE2Q�R���K� B���Jɛ�̱e �?�V(�%�'�
!8ب�$tB�oʊ�����}���ɢ6:�������}=�b�Z���j\D1p�9ߊ*���<��Ӟ�Uރ�1T}�`Z�T��.�:����u�o
_��l����)�JQs�{J`���Lu@HN�]�/����(e!xhj�M���dOG�=]x�K�ӧe��mv�L�=$�+b���r
2���������Sg�!�ut�V����<��=MNY]'�֭ C^��(�
 �,��&��B�ҏ^+�	J��P�qM[&��L\�%7�/"��I4�X��"�z�5DE�8[��xD���\|�l�v�Acĝ��נ�\v�1�v.8B]�rĂt�6H
��g�
v�g�l�!D����!2�᥁8�������\=�i0����鼂,���*��Z>;�G"�M���BQzMP���� �[j�Q�^9	�;��t������x�B�NqC�N�UiW����A�;f� �L���d�����K ����.�T�K���u�
\h��g(���X����w˕-�e�?Wq!eؙ8&��3��+��_�U-g��ļ���dˠ 0�\�'Q/EV�u	��	p�r��8��,>�S܉��:�`pv�0z���!l�6ŇL��kWbq�d�7�
�!��E'XEmS0��n� �^#�ؠ�ɂ�٣�KN��mc��sdI�A�������"һ7�
*�iĸN��̧�$�v{��� ���su�d1����A"�J����&�M��A|db�rh1�F��/+���Q�/Kt�#�l�PFͮ����}2K�'e�n���&�»w�JkѠk^��J���ҿ�6�H�g��#u���Ƿn���$(��e�}�`f�*R�ơM)f�hm�
2	�~^��t�:��u��*��r�"��:d�t���^7w��-����>=�Xqt1a¯�,�u����<� w� ���su�� ���($OM�V[�Z�ظ.A�e����Y�:�.�c%���P��wdx��#��!x�@U����˓�_�Gʚ9M�L��jj�.�� f��_R���Ź�]��8��t^� ���1�C&��4ɾaB�aY_�C�i-�Y����:FNS�Z�
���g��`�4��\,��Z89�ė��qK�?\�|������~QՋH	2����{v���_II`uQ#S&%���{�D�~�!�7�v��b��J_����ݩ������n�O�%�@�4b�6��k�j.j�͓�~�mb.4�jh&���B�nK����#�;@ke�0[���2��!4�;��
U20��R\-\�g;ˣ�O1r+�ً�?ۖ��ۮ{�p���L�1���"�8?�}'z?m:�CZ�wҪ�xG�؍Iy�<bz�A��=��Mjv߃:>]i�I\����v`��
�B�{MckzT>ا����|U�66d�AO}��� ջ�#>Hx�;�c��D�s�1Uo2��y҇L���&@W�X����l���i�@������<�%���ٵ]&��WY��S�I#��y,2��xNP���ҹ�3���t��`�-�/�N!�'V�Ә��һ�&�\jt�-�`���f�&���ΐ%���/���<8�g�#m���wF&���o�,���m@s*�#�Ӡ]��A1� �"͕Q�7K7��;9	j8I�6+����)�I�.�B����y�$4��z.|�>h��ƠW�]���\�y���yB�d5��q��e��$X��%�Ca��\�p_:�u	̢V�R'ݗ�Am``T=H�lt� 8�[�AtS��6��e�y�:��l$݆>�c�3��i8�K�mͻ��7N�2g�(�il_B�(��4pħ��s��P�hw�E[��8��/0'(^MS��By��l[f��i#����W��-$.�#2��u��F�O0<,�c��(�f|�+�ggߎ�o���;[rĶ�s"�j�DJwڶ$�ԑX���uD�g�F�)��/����,��׹�����5�0V�p*Qm��uSp�d�p��*���&mh��C��R�,>�N* 	i�� 1���r��s���/�3%B�b)�b1>ln9-�KM�S�2���z}�W��f$���f�Ma⟄mϓr���$��{>K�����e�q�|���B'�.gk.�W޽�W���J���'�V�ɗ�z��* �1�V�bqll��B���z3aB���Wl M.=a
���vs$�EA��Ť�h��k�#��S)�6���6���w��)�}X�;��ͪ�Ei��0�,�x���,eR����BhT����ӓ[�2n�=y/0�<��iYɦ��4��(��B��[q�>��4Ź��aT�����_\�Kx�*�>�K��)��Ӽ������:ee��Kz%����-�a�D�����NDf��v8U��AD1�6�8��49y�W�^�Èy_yW%����ﶎ������䩯���^�g��B�v3����~̜��C�$�㺒qO�QK����� HV(,�~�"�������`�@����F, &�I�1��0`?�Y�=�����b7~���6}�z�VZB�@�a�2��������2�����iɑ:�V�� �P[=.�N�@U�4+���).l��FD�k PF�'��c�'I��xD?"�:jL�tEUV���\��ieDټoF_�q���x��
R�i��[��#"��Fv��(�oc9��p�֘´0��'':��tצ�uw�J���㯈ډ�u�
^%��^m�T��:ǹ�O(�M��ʭ�m�~$.��;����]����Au�#��l����?p;���0�{�0�H�@mڷek��a`JH=bERƍ; ���ϵ��^��K�r=��6i��?��&�Wn�]$�Y�M~/���Z˓�ЊD�YN��xJ7�m4�oF�"M�Ș�F�E�
"�޽�w3ıʵ=1�g6��������(g��}F�&X6Z�,����?�%]�!d�|� ��R������2��r�%��p��
��ٳ���4�y��/�pi�Ty�j��$c�:�*�8��sO���^�M9�QM�Ϙ���b�����|a�-��
R���XFg���O���yfL��R�x:�qE��G@��rCX���r�eW�V�������%v���D��������Gpγ�~��N�ķ��ҡ�Oz�Ne���%�{�7�HO���إ�|�Y�rw�@荗%�����釕���eZ��0���ޥ����a�+�Z�OƠ2p�O��.�N�A�b��5*� a	V��4#Ghvg��?�j��
���.L
�9�!����"�L��	׻3R����uk]���oSLu�~��[��.��WD�ľ{|]\���>f������u�U�V� �w��S��QPM^V8z���I`�{��>�"��Ӏ�cg{էE6�P"<���Bd�{��hm�}�t�_ۋ������&vl�1+7�#_u�]���e��]&M��8���S9@���!�e�:�Cv>�]�X�g���E�'�~_y�U��E,�3���җ:C��[�������в/�KB �EH�SB�ј���&]��'���Ú��ڞ��`탯L�\2�Ͽ�,/Y�+�{�	���E�s�/����i��ҿ�Ԭ;G�����b'��499dZ�����
��{���s�p�l�$1��p�e�K��
'��.�ME*˓Mޕ|b���LT�s'���<���mu�D��������BW�p1��F��Ksx9�
v'�gF:�qv>��K��3	���$�W���/�����A�È�˘ƒ���.BҚ�<�� @�}�>v�t2�<#�_9�_c��V��Ņ�������d&�Q��r����d����f�N�j����A�T�h-}{Q{q�g���k��h$b�X���Z_��3��Àec�	>s�<~w�l���Y������T�k���I5?L$X��Um��گ7�(�M��vz�+��̧pH����.0���]][+׋�v��}H!��.��$�?;a_$WL������ɍ�^3�����@Z�e-�n�p���a�S���i�#?4Xv��rQ����L���k�;���y{��G�!|R�#p�dJ~��}'��m��WtE��%xYF,���.��d��^���⋆($�,Х�ş�Z�ףo����N���~|V�}cs/��E�tS�_�G㪎��ŵ�/�ak��GO�A�]��6��M��%����O�
�V�e�_�X=��S�,)���
��Ǫlx;�2��!�Z�K��Nވ��'��?�G�����B�	�,�N����i?5�.x�#�Ng�����Bh� �7���Ҍ��q�]�LT���yOKw�/.�㮈)�ᴅ�vV���8��6�4� ��{hU��h�c����-����y~�D73Fθ�AU �M*�Uootv.|Yn���b�Q�Q��<C؏�,>�^Ό��EBI��1�a���	WfW�(:<0غ������p���5�4k���G�~oS���zZ�	J�yRݭp��(M�E�������,Z��%��K�-��T��(��>{���'�_f-�a�2 #�>e�J���ܝ_���C���C�F�;6�vaܒ�Ȁ�c������e���τ�+��B�e�j�(�TI'���%1;�J�?��<�2��w����<�t]�杂<���e�>�k�f@������Yxqt��iI$��T���Lؾ�qv��N��U��l�軭i�>ϭt�G��n���J+6��|;�>�]�3ءZQ�IX/�K��^@��fGrt���3K	G)t��w:n]����?�ƒ��FS�1�e8<�5%T a�������ݣ2�sb��o�TT>�E;>6���E�,in�7Iq���{�<F�⌑�l��`z�Qº��h���K1y^r����ܯ@���8���I-|]Ս�5B/���ߧ��ˠ�q�dK���^�GwC Ҫ���	�Y�o7R�r��������PFy�+��g��i֍�3����"�-n+�F��@i��W�YWZm���;���%wL�V���"�ܼi�H��n�ц��גE���L���<1�Ц�l�ߘh"�G����$�(9bKzPˊ��9S�3��p�Nq��J �Uy���|�	���G�8�{=�Y�E�W�m��t#�U8��׵Di��Аյ�V�_�Fl�����pԫ�I���!����ǃ�2lTkS[&������E���sG.|M%�ۺ�".�+����;�ؼ���Ҵ�]��w�=
���	/� d�C��K�f���b8�{�R{�)Q^� �V�K�=lE���P U�l@}�kA��� F�ɏ���h�>�tumgw�ט�Be����dm�����ڛ��1H���,#	�?��%�� �c]��>���Ɂ��I��5�e�(�֟�����m�����l5���aj�i<�t5,'R�w��KŒ:x�-�P�_��+vܯT�U��Q�'i}�zl��	�B�N~	�MWSӻ�"�"�#΄��1U����+�Y+����0%�d���|"v�Ҧ��g��+�7T� ��Ñ[(e�i��NK�1���.�U�����ySz{Y�' T��I2.=�Y��N�y��5��|�{h�s�Ai�|/�r�B�妸��}К*��Z@i-}gD}�����g4��Չ�:��{�Ĵ��P���
���F�����'A�/>�%����K���|�W�/g���Ǐ�0��6������5����S�8��b(��'���aq�@K�a1�� �&v^�2�JrFіbǂ��=�K֞��N`����$��p�kr���}�M����a?�8�J]�v!Hp����
|�?��{0��eD�8�T�'�����.+ *&�Wd�d��eBFcs����w2�;����,a��G��80N�%��E`����e�;�#+�ݰsaj�x�<�!�zU�b߳� ɛEX��c�����=�\���YY|���w�E�:�p/3�ө�!�_t���y$�lF(ͬ!�'�j��)ܵ������1ܸ���2p�I�?A]�7v���ý�Ρ%[D�?��?'z�F�}�ʞ�ʳ��?�#B@�����!�4��7%�� ����P�_ֶ��+�(y-n�\o>�?@�����n"^�p����\�l��Π:��i��$(,�b*�,';[I��N�g.�YP�2��f� �u��4�X��,�{���?^�P�DS�^�p�B��+C[AT�+b���f�"��7����>����s����s���L&�Z�й���O�uk#��7�*�>S�qxhe1�Za^�����n�w����<�b69uVA�3c��^�wS�>�'e���\神��9T��V��]w�ނ�'��:gW�XXJ��������V����='7ʎݪ푅"e��]O0lTl�A���鴣�
(�l�;:�	+4q�e�����"���C�J~fz!d�6�h�L�ҋ��UG?��Ѓ ���r����Ztix���>E�yT>j
���O����MQh�Z�A�9��a�"./�����?&�
��7Y��H��������P������[����˷ZW����y�"�<��ZՀ�Ͼ՝>K�ם�҉9���8�s��@uW1�/,�t��8 @>�k�?����9&�r��x}�a��C7]z�7���DI-eo�Aҁ
�IZ�G��֎!z�x�'�SB�"����5�!�䤭p��&"�&��x܉��o�gQB��nѹ�^�c�Dd:#m�J{����Pm�#T4��Ŵ�y�}�'Ƅ��d�F�s�P�$մ��
�y����J��W�ꎅ�Y�8�Ƴ�=~y0il�d�`�mi|�Y`�� �����K�>�`�.��C��<��i�~�W��OG�HY͂B�_*&R;�`�cL��nU�}�2��ݼ�YX!z���B?�C��^4j�� �螠�/��vt;߿��/{�H�C������"�c�~��:����S�����M��e�aJ��:��s��>7�|7q­���W��GVC��g����;������O�AU��8�+��4������vE V��s�6d�O������<�K686WS����Pd#[���n�m�K@;KD<I�=����Ԍ%C3֓��J��T�ػʌy�msa+���O�!� Eo�B�;��tX�N�vK��jp7����fO�.���_���#$�p�&�kac�dG���g1\�&���Yp�JÌ&��tO���J�K�5�������~�1��9��]�����;�� '�U�{�KΣW�L�Q�WY�Kfw#�����)>�ɳ&N)��'O]����oaڮ�������=��B)�M�57ͼ���P��4r�6
.AV<{�C�����0��S;Ŝ]�@ċ��l;׳ܔ�Ǭ^��9%�g�����[ %8\�Aj�:>f�8�(�n�6 �� $��,�>��f��k+��1��Hx˛���Μ9}�߀�Cb��4��c�R��g��|U���=�Zu��d��R꫞���H.Ӎ��;��	�z�q�ۜmy��2^��XF�����C�%�SM�*�~�w��C��X|�3�M��3M�=G�R	��$~� <���7p�%�{0o��2guz���\���|�1O��@�^�W���0&������~;���.U��j����Kz���1���ib;��R��	��%��8K���]�X� �)�_��MQz#����ąDda���z|='D��v!H���dY�����%R���l��*1"�5�J	��#�"j�ק�-[b��GD}����9�*t�DW(�&~E�L�'�O��.����%�\�9�d�8�5��42�>
#q����
�h�[pg�v-ܝG���ܕg�Z�h/~%Ǣ,����Z`�Gt�mo���
KP�h6�<w���p�U��6�f�X��|eؔm�J͛_���m�{Z@V@TL�4��@v����n���2g�G�`�XZ�U�L�u*��k���|�����>q��e��r���>k�w�*���e|	�>�g�$�g�]H3�;B��fYԞ��/z��w�}���J�Q�q����юcW��"&ﵫ�ß�t,N�Յ�H��0�$����`����E��I}h�I:F�j��$ߎ�
�&�ț(R������<o�'_([d47��*Y����d@ng�(�3��
�b�����Ap�C������i��a���g������� �c32�^$2U��m& ��I�s�]��;��b)f���ȟQ��V�.��'�	�N�$&p>ɉؖ� hv�y-K"�ii�%��XJ �Kױ �k���B!�e ��.H=�ȁ�~&4J��>������`=0�뷈 o��W����?�T�Z��(�D�S���Ҳ�)�A�7��˒�������YܤimV\���"�q�J�'��}9RW�����q����@ �`��K9�3v}��i'W�ģţ���$�6�ݮ�aQ�Br[���A�����I��S��H���!!�!`��"gz/B��(��zUo�X��$�sLC}�N��z�z�U�GeK0�������r	W�x)L�c���A8�������k�El?F9{�.�c-�?Zg~$Ğ�8�g������7ג���׽Af�Im���:`����Jm��"`��*�~��|�G'/S�5�!�a%��6O���/]zT��裛ĸ�Gr�����"��X����k~D.J����UԬ�U@
̊t�pA�Ԣ;@��kFP���C<�{E�����j@�������`f_(�IP�j�]QHG�n�m3��P%)�I�1o�cQ�6�C��q���9�Q2�6��=�J����e2�T���9�Y�<���טة@@�FK�T�%��4�ZO4�?XT1�ce�CΖl���~�=����
7B��{u��5��鶘NSz�Y�����d�2�^S����t_����:Xu+�ev)%�_����7��h/����ٝ��\]H8�9SE�v�(=�/Vn������� ���l�T�����$��|��Q6�Ǻ_�$S�k�2UX{o�l���z%���Au� Ἶ��M��虼#���Ә6��d/��*X"�l�A�0��}�iYN��d�pޒ��e]+� TS#أ��Ӆ� ���BN� ����)~�[�I"��<#��]3Q�.s=q���@���*%So����9�����������-k��$��C�������A��s�zZ%| ͏�^�p��`���ƕ�o�� 	ɦ$cЬ��&����v�؎���g���Т�/�M���練��l$H��x�+�l�S�X�e��'Vig���=V|߷���}�������2q�{)����� c�e�m�`��E;y8�֥Ab����%��lh�oe����K����4��,��)@�o�;��e�iF��k�� ����<�6�n^b�pׅ�8:z{5l�Z��4J:7�=Sѵ4t
:�Ҝ�0��C���Idߚ��E��4�98��rs�������FL�k�yE��zL���t�D]�qE?4N��܃�Ʋ�j��3g�<�i�G�7 [��pj���³����(�����/�@:���yӠ�,�5�&G�¤K�A�#T����"��2.���U�UK���K�Ѻ_�������@`+�V���	��?�F�ߞ�g���B��5�	�K�;K?~L�*A¦ea�K��<l/x6�ɢi�.�.�f����݆�8@$S���?>���GE���j�����W�a	��jU��((�㿵��'i�܃V�S���P��L���M�\���xaJ��U�K���k�$�1�����)��G�:����Qv�t활�	Y~��1����^���|�B!���"�;�������	?��Ƿ�΀W�����fJ�Tm͌�3Pށ�7I�P����K��6u�x���t�f%&�R�K�q����Ъ��X��!X����Rdu�^�[^��q,�@v=�V������Ɣ�!�|�Ar��{���{��[̎����Og�7��5��<�xԱ�]�-6���>A��U5��^�RG!��$�u6����r>6k�����;�k�F�Yj���yW�/��ڧw��
p����h�=�4�1��d�lXF>��nԬ����;k�j�5���m�%�z� ���Jq^�d�u�u���)E�bJ�o_{�j8� th7J�e�I+��i`�.K�Њ� ��|��FD���(5�m�Y۱Q��S`�5�F�4�� ����%�ɡ2$ѓ'�gp��~,#KH.r��=h�L��$�V6���B&�sߧ���K�<a�[I�6�Ҡo����h^,�b&0>�ӏr�D�vc7D������y.��p��]7���]v^RM��?�I���Q&N%F���c�Vu�`f*���	�n�Ѣn���u��n�!�5~����{O�27r��Ug�C�gM8Q=?��t�B�up�|������Ѭ4�}�T�腖V��pV7���~���[Ň�WI*�7Y`��#M�'�B����'ͣm��r��k$�M�W��b��'ʢŞ�	�A	�R�]��۔~yP�b|�!u�m�� G��3��Dګo��-4��YuӢ��2/�� ��2�����M�W"�8
�^r�}B����l#a�\;_`����3U���1s�{C�M�D��xތ10������P9��#���pb&�� ����pf�K������AF��o`Ȼ@a K.T=�7�C�/���o��
ʮ��7�7D̨�_^E$�U;�Zs=�}�Co�Ҝ���z�o:�R������q�	��Z��Y�D
�WbM���f���q_a��q��H��K�eP��N�A3|L�����d�4.8��:�ߵ�FIy^�������b�KL��;?-DrD�,ӓ�I&щ���^�֪LE����8'�z�����hg�ؖ��]�R�f�}W�<��yU���}�B���Eb�w�B����{T16v�Y%�8K#�k�r�A I\���0ｵ����EX�OJ]Cuw=��Yx�ӂ`zDH��R��Km�����?���^�����4�����e����v;������/���5ث�^ t�h����ț��b ��P�I����3�l��̛B4$����a�ʕP�Ӛ�k��:��8��0���h�����b���׍�b��Y"ZE
/�_M6VK -�I�3DO;�c���Q�|��#̬V��n�QF��S��|��7�0��,T8N��O;�C���a2�d��+f7�o��"�}*/��Br	��ay:Q�~ƌ��k��d��A-�P�׎|�pTb�=�X���i�lQ}ޥ/���nDɂx�'�s�&F.�����B�9�%\��{��3E�6���3�,�hQXƴ�94���NgV��/�n��ϯ�n��~A;CtW~6U5x�	e���� U�e��4��H��#|���E�����f��@hi3gD�Y�GYmT��H�.����2*7�L7wY��Y�U�g�5���E"��`.����8)�7�Q�Gf 3oYUޙ�� 9��׃¼Ą���u9�c�h�r_���vԤ�i��z�'�Y����菕��Z/��G^r���&��ڑ�<}mQeM���~��|�m�̣��O��w�ǊM5�N��1�3�(r����qH����q[&�ݘ��>p�Gv|m�̘�~�'ޠD���H��SWoE7(���,���bb��I�:n!+��$�fs���rY�R��R�ђ)U��6\�Ay,ote��lX�,�.��
h��@0x1���np��?6R%���e�.��U@r\�q�:�k�6߼���|]B��b�h�L4�6U%o�dl��fR�Y��OΑ��.h�ć� y��Ӻֆ���e��n�,[K�~�x�HE�l�(��]��"���|�~�fx�'@��{諵]kݻ1(��P�26�j��ڔy��
���ϸ
W���,��߰���w�aR���<�c��dqf)�oɈ�{����9��T��Wu�J3�:]Y�S� ��"K���x�����i�.��UH;>��p���{�o�$_�p2�|Mť_�S�Lw��2gD�}�{8�@˷�fTE��[�B�2LM���Df��У�c�\}�9Z�]43���NI�q4�*^�%��h]��۲邮��\U��ZL��1/w�V�X*�5��rr�`����Yy8����\g!��/��v^�LB!�g��(Թ�9�+�W�Qg�6��~U�����'�ʥO�y'��ǋ�F���}	� @�M�R%��Gi��zH؆��L�3�n����󊏿�=�ɁK�m��������q]����aʦ���j���q5Z�f��J�f�� ե���Rk&]Y��i�fM1>�M�8���x|@������6QR�i�	�U�(c�<���"7�̬^�u`� ����'jWm��&hh��so���� �|�Ik�N֯i���V�y4|B�4G/�\��r|Q%-;�Hr餵�+��Yۡ�%U��YvN����i�e;�X�N��v�|���-�)�ioMĴF���o��W�l��P�^��<����x]�֐��	Qh/$I�@��#��
�I6����-�ۆ�1uZaա�������x�y�Cm���>�[�rH�3\Z�1�0	��#B`F��ѵ���b3�>㯐 ��0V����e�������a���(��(@kH�@�=�	�ba�gBr�z�6�q��H���vr�V��,��'Yу0�7��Eň��Y�tT~���J���J�+W��59�,RIU�!R��vQƦe �G��p�m�T�un��Z�"����o��vW�مAҋ��%���S|:�����O�Q3�W�
�'UU��aY};x�ώ�%%����^QTOQ������r,�҆8;<�R|y����kݎge�%ªz��4�.#���?-������!��N�y�R�đj	�����6��8�_^�kD����:�u��c?���4�HS�wdZ}����m8!�K�\����@�f��쎝��t�bE�������[m����I>�:�1�o��(L����uGw������6�"Tƀ�A�SM�?�c�{EG�z��{��ww�6lb��2�)#�"�}�#�w��dZ�<��6��
Ze���%-�JR����m
��g���ǌ{l(���@���|\MA
C��q�(3�� t=;��V��B$�f�?�Ի�YAx�QY��$��^��N|(����K,���Y�0��rE�֝���=ك(q��37��!�@�x�����&6vM�W�{�|���X�i "&�X���}�3��d��K�R�=���i�2�ʁ��g\��"<ķ+RM�V�3"0ؽnas�[$$��Q�,.v9��Bj1�\���耜�Bh��Go5�il��`���O��UI�(Ğt����a�U�3��u��n^`�倿�!�^"�x#�ސ�K��C�;�M�d��Y J�x��p���ؓ�@��ԡ���}a[���Z�B�����d%������ĵ�F*�:���u~�5�.&a�௎�x]��3�ѦR1�������o�
�bAq14l��p����V0ic)�I�P1
�:�<�HhLa��[	TM��l3���X	?I�h�N�B
fw8ξ�ޛH�N�����?(�[[X��V�&��Ě���/�q���}#����z�GW"�7���B6(.����`��3����\
=�c����M�@�����E��S���i��;��-�M\�bs�s��b������;��`qi�H�\ZW-��q�[^�M.���V��!h�H����=؁oc�ͲlB�Ǟ ���YFt��k~s"�|�����:V!��}����^|�j�Lݥ��& ��uw����@{�}�I��p`�'g��z�6�\�>��8��n v��o����qU^����Dt2� ,�LVX�|�*_�.�a1�ޣ�˰��#���[S20u��7�8�>�_�Z��P�L����gn,�/#K�ƌ�͙oFښ*8n"��;�+��r�
׏dpL/��	���9��Wѳ��	�u�=���{h:,���� c�x�������0�>l`wx(���2����=*��� ���wn!i{ѩ����i�e*���"���!��JN��V���r���x��!��q����!�8%P��s�@�y�$�H�K�nHGX�N�v�<>%�3�-�As��*�cy����w�FQ�Pwq���{<�dz�������C�HǘK���$�M�Z6���t��7�0�@Ff�A0��i��<��W�?���8ؽ��F��b�D����E�o�X� �V?=�G����9w�z��\3�8�	���}������j�9�wygH��j��)�yw�#�1ƋW39̄�k���P��M`U� m(~ �3Fσ֧^���o^��a�!�O��~����g/��a�gB���칷���n��|!�[��9q.b��J'w�JtՃ3�5�n�i������/"E���w�uDڢ����G��ɐ��:g�D�A(:9*a0;�'���#�V�N�-Y ��O�*�nD�t���p��O�;HSGb�)�6����ט�<,�U�&�te�Wp��u��C�fV?o����稓��H��VPp>���%g���r5�'�:El���~@���@��}.<>�K�$|n8�A�%�yt�@!�j���&-^o(7B.�^~��n�w�pW�i��H�!�\o-G�0FGv ��߸�c�[^X��v9b�P�w�>��WL���.���iP���\�,�.�n5.��FɃigrT_�<ω�N���e`�>A����1uB�ܗi��@Q6�SoT��k��gYUQ����$����� ���iU����9���V��2�E|o�>w&���,��B�%Gή.u�	c�!��gB�6���l��Njb��>K�>gZzZ=I� �>�H�_h�:- �0�@̏paS�Q7���SS�+�4J�>�e�z��z��dg�$5�w1 tY{],��_�� ���H��2\Ӆ���],��V��B��� ��*�Z(�"b����Y�K�Qx���X��jt�+�3�)��z�����?~%x��1�ơ��I�����Q|���:�L����i/;��{��o@t��Zf�lEq����i��!l����7��6[Ǌ:F�*C/I�u�Ճ $6���:�7��Ӷ��j��i6�TY*{�+��F�k�Sa��H����?̗��EO�&����n[�COܧ�s2zU������z�[=��Y[z��Kh���L��-�b���ڜ����n
A�00�"���|�Pa�r��j��}y��N�>a���C����W��YJa��\�N��iCc�M{`�@��N�@�����f�
E�$�G �p�{,��� 1�yKn�K}Pᛜ��!�5'�h�%Y�/ !n��ᘀ<>�SPrQ��VCV6�����@�wݘU�Q|�%l��g��ݛ�t�oKm55�<�&I��ڞݚS��/M��:�{��+�N�Q��I��^������)s#�P��pْ��]��♄���Rp۳H3��ϟ2nJ��%�`�Z@���.P���=���:`�e'효c���<�؝��Q����7��=+sSu�_H��������5�w��NՃ4;:�)`�Wݔ�Hְ(� ׅ(�m���IUY�b�N8�<6�^Z� � ��US�3z�l�zǾ^��-�ѕE�K�Bʑ�m �
$�Vm�&�q4v{����6k�N�L�z�����)$���ޣ^��V�Ot�r���t�M�q��CӠ����H�h��G�"&ho��>GRoDض�&�'`��mU,�Vݷ�rGt��xF���J�Đ��,����c�-&��gEY@��/=U�+�1�y��K���ӀN4��fuUgUؼ\ڥLW.	�<��m校t��3�e�bj�U�2φS�a3g��0B|��${y�I&��l�o(i{r�j�J�/���v��Z�pK�kq�l35���������Bq��;ЙGB�-�ө�ʌ�@���E��+8�Ilv ��߿��F�x���q8�<�1��+��B2Cz�B�������u�n&�T#P�FT�-�Z��D���Ӝ7l�$���C�@5[3H��|�����0�]E{w`���0P���?	��m��Ƨ���p*E�Ǧ��E���R
�b�.9���O�T�~��6w����.L�%�g 9k_ON��#"����>����*P�A^W�?vz_;�e���N�S�����;wp�FP�x����F�m'K��ٛj0�{؟D�!��2{G�T�z~�O��qϸ:KY}�`�r2��ќ̨s�KFps�~�`1��MZ�3K���r�MPQv������"�r�85XuMg����s?�=��I�Ć�O�w��]`6�%+���z�)s�����Z{F��!n��͐������V �=�$����q��N��яC�6�{���E"^��{�y�S�A�&��w��g �|��<��������@�)�v��0��3�@5�f��X��_^��uQ�0�O�)��#m�34�����e��ȍ��·��Y��e d��{����z,���6�~�4459�k_c͆�v�3`��gi��xi�n�v�6��yJz:�y�5x�n�7	�0�����>o��B��A��(�r�w|���{����;���×���
R���m"\�q�4��z9O��NzN)e�:��r �L��RK���%��+�iyZ�8�͸oh�I��qh��@h�<v�kt�^��M�Qv��� ���!<2� S[��}��g[�qW���<iS��~�[Jr)�|���]��mJ}�l[���K�� �-O�	ڔ���f�>FjE�{v�m� �f�c>� 6���� bB(�����x�F�&������L<Q�0���f%g&���\g�l��S��Ha�s��(-�o���nL�T�~P�H�2��$���U�"�j������M�ٜ���Ԙ�#��<�k��{���W)�e�C{|�P���)c.��p}f����V����2������]fn�Ihw�Bb[�F�j=��tFu�I`j][����>!�>��^Vi�x�0�+ţ���ė>�rI�[�c��ź���Ĭߦ��r�ו"-�Y*3q������!�7�� ��m�HmP�/��t,���2;��2�k�{	�:�a�9~�:��St����K�\�a���������9'{R�YV?&[z7M�s@$B�ې1*�f��玴��G`O�t
-FH#4�y��V�~6����`�f��m:��_���9��o#�E�y��2��zü:-��=�i�ys��vn�l�v�MX)�P�š�F���ր�d?I�~��m����.1G`��ݦ���%���,�=ij�����n�8뀮��I`��|�$à�S���=zU7�7�,�t�8b�\	������l���wN#���ބv�:[7�*T�kA�_��X�-�LD!�B��~��`^�;��*�<!�j��I=�gs��-X��A�������nc�
�P��hʲ��j	�!=w'�>�n��r�J�H�R���٘�XhSJ��C���F/�~��[ z�q5�Cm`E��5���LWMJ����7�7���_Eb�@��	�bnzkg�k�o�+���k�����}v�7=qh{��-<I�C߆�M�����7M10�!�ڼ}l����r�v�}׉��e�a�[TE��z�0��sLK#*�&�.����28p����h$���;<ew���}0�Nх �N�Yg`��h7�J��l���E_�%4#k�0�jS�䘫�f�I�U\��"E{��&5�3�!�5%�9�_41]X��ܹ��f|�q6��d�k&�URK�������}�Xk�Ӭ�ѲЋ������k��K��jY͎�BD	2n����̂$�����]���"uS�3
�G,�����3���<�D���)�_!�����
�;�Ȗ'�T$<ͯ`��(���&>������B&��r�����r��ܬ�f6�T�5�T�A4�:�9y�0����M�F� ��l?��5��JЦ���P��ֱ��߆чe���ԝ����F�d)�h��Bn�����+�-ٸ/S��ϔ��6���x]�c061��R�9��V���`��%�a�B�[~���A�q�G���E(��-K4=��P�Uk?7�q�r 8��`I��Sd,S@:����MJ-T|3w�I)3�d�0z���$��]�2�f�Q<1���F��v ��#��V�D2!ק��0�Ь���E�Lt�I��QZ8Z�@`��(� ����i��S��~����\~T�-�=�4�Y��~���
��(p;���P���n����aͩ��*�6˶r����+V�}��������}�_�I ��W�MU��ǃ�> 5�]#���7i�NJ�8�N�� �`���p�~k@~J0g[��I��I�E��l���UV��>Ӿ��&EM�m���J�Rt㢖��B���N� '�൤Ip<�����Gyz��B<r
�޷��W * �lL����0�����f��)�8�B<%�Wk������d���Ϳ�{� 	b��&�l�*�7����ri&�6y��>�5sE�e�޵��X���t[To���i8�J��9s*�ǟ�g�SKq[f2��t����1�R�<	�]ȱ����RI��z��>\�����#�=�9�{��ކS]�1Vw�=o��Rq�y~����V��4�a0�';k�K=�:88D�O'���Fj�Y�M�нU�qX�k1���d9��ܮCf�/D��4C�#�^���Oh5����0��N2���?�x��3!k�;�D<��=$�4�q餐.�kގ�)���yAbz���a��P�J_N�Z�!�n�SmH'��:=q���������"m��5����w��3�$i�v��H��8�7�~�&��r��ѽ����d���ҿ����֏AY��z��(��]�y\�_6�!��;i������m����De�[�y�^��Jm�Y�̗�n8y�A	6�I6�̓���g�\�([.tf8K��'�'H|g�k��\�����7�u���fC��!s��b4��f��ȓ8���xa��o@�m2D����]'{�&	
ل_QwG���Ԃ"�S�����+��,� t����#���Y�
b���-�Jm k�˙��{J���w��z:����<I�f�ՂxT��\���,7��0�]~��k�jֿ�	��ⲙ�]�F[)
=SvM!��c��뢭E"G[|�C���2��u2��r#Y�&�[��WV�O8;\F�%�F����׃mN%���Q�z�.�/w���٭��C脌#�U����r�\��ad����H|��O�)d1 ~�p�rS
5)X$YWtNP��pos�U\�����C�b./�a�
��6BZ�;��R���j�̎�m�	a�疒ŒD#�'��(��+����7`Y������7���1,���̵����kL$,��3�hȷ{l���ڥ?�*�8�[f��/��k�����r��mTMI�K T�0~�͇�e�D������4.��i�iwU�H�V�N�l� bV)�Ï�OLxۀ��3�{C�r��8������..	����iu���R�OY�M�T �(͋zG�l_)�m�����{Al)�:�tK���rН4�����5�xkl۶e�
X�~d��Rڽ�S����&�h����E-PKLmyj���Q�lA�T�csmU��@LO��H7(�u(,���evy	�h
[�HX���/AMO���T1A��i0RPV�?8�
G��#���BR��ֶ��t`��ջ
Zs�Z��v��@@��}Ĉ�N�����cD&_%��VJ��^�D%�U��E�=�
yn��H"�S�q��pL���<*?@��q�Yk�����(fxoW�����٬�����wH`og7�O�����9�r8�O�$D����������35(CO W���=�5�ȶʀ���a8m��N���8%'t?��*��X�F�����S`����u�6R
�b�s��25�b�x]8�%��� ��%w�t']zץ����q��|�+øm~��������2ڽ���cp�O��P�U�I�� pA�W�y6R�D����{s���]��q�դ/�.!V��\�҈�~!��V0�TQT�Cy������遫�v0�
�_�#U>�V��vO(tw�<��à<�}?j��F(|����v wo���p�Lبbʄ�+���
�VW����������h�;�ÿv��!HF8*��	'���D\���7�8x�z���䋞(F9)����٠���S�X�\��GF�}T���J��~����Q���u�3�U�L�5�]���a%��p�+#�x�f�H�U���A��xl����.ot;�� <�Y��-Cʫ�wL��S[[�B���YJҸy���-C~���J�|#J��;}Ͳ;^ho�r��Ģ�$��rz����Q��T��b�e�:m��
�F�$9a_w�'k���;�����6�����䊦����F�l�N0���%�m��/qJ�����2��P5p1a_?5�[���{!�Z�?�������px��$�GFue�����'�۽ͪRx����A���|ƻ�)���h1V�`苴�K
H^Mi�v�-�*���^����������<+TԿ;wy�<Ԕ�}r�oz�%z[�t8~��{/GAj&�*���ݻY���w	i�Q�MaU�gF��Y���.G�8څ�+^���i�\���@�n1�٬���������>��-�>@,#㻀���gO��NXH'��4ޞ�L�!�D}���Ic]�؞��V�e���inP�6��)%�@J{9$0����1�iuB��I�E�m�d�"����$��z]3��ç�M�II�c)CiD�'h��ۻ^�݄�z���wV�P���<��T~�g	�e��}��|�Ёm�rC����!�?�Y���Br�t�Sߣ>�B���vu��=��Z�oh���=�ݐ�'�	���R�3��=ɻ� ��"���?P��+��F#o�$��A֑N�xB:�֨R���+�ڂ|+a��X��N����uc��r�o-Lovg}?��J�s��t�$���k��(��gp?�,ʧOUFf_"y��b�F���S���Z�/U��Q�C��+��_�$�M}%�*�͚�����
0,�<����7�lW��R�-^v�|�d'mܧ4^4vt\���8�زq�1�&UP�5���n����E��4|L�t�Qπxpm>}r��m!q���І=�����>��:�VS�,.�\dj��J-�Y�^ҽ����;3+Nd�#|�
�9����,�v��$�({3�Z\l��O���#��(]B���~���]C���3Qh��yГ�W����9.)�/�.��z_���/�%6婼�P �lݘE��D�\�J��YB�Gǡ)0>iFhg��{�A�8m,"N��A����4M��t8��� �>Q���� x&�(��c� Oq��V	M���u��)D?K��{�XG?<C���ľ�Y�}Z�y�`E�O�
��{eeW��6��
�DMHhbD�rXh^�L21yu�5dJ�S3iͰ�0�U/@������P��&:�K�0�K!/Uiʛ�9�F��)񄰓6�l��Z&P�d0F�+(�~��Rs���� ����e������e��'؊r8�%9�%Q;+�eU����/\�r,��`� �&c6:���MN�?[p)F*�1t'p�si �t�GP�#��Y�������G��A2[Ȉ4����v/�;��{t4�o)����*H��E�i���^�Z��&iq]a�E�����棂jϞ~(��tB����?�L�Iu��뾏��r����O6,g6e���k�����Hi�������1�U:+�
�ƛ����5$���{���j��� ���/il �G�� XU/JTu�2�̒�tS@]u��~)�^�\l0�c���`˽$��i2U��<\Q`��$$d�e�����6	�N4���-��Y^(�?�#s>cW�uN��U�ۃ?�*?���w�-Z�L7�8a`1�xȥWt�ҫ��J��zj�b(ݚ,N�|�ό��m��}h��_Ə(��{��O9}��VϪ�惻��hMv<g�s�7>C� P�w5��g���[_kx�I�R��)?�.�qh�Tz��;�x �Yu���� F�ÖB������}әh�L;ּ-��Ӑ�G�LR_���w�uXy�2��ģ��!�0/�3�ic�X��+�(8F�x.	����0Y��RGa_9�t�+�{�S����N?�4��e�)m���Pv�aЙHqRA�@�u\���'
���`0&� Z�Js"��s����W��B�9�7��8���Z���vi��T�C�c�g�����a]/���f�=���Ȏn:�r6DqZ�EDMI��a���cl���Ng{B��>�[߁��SV����ݯ���w�q��z<'<e5�^ʹ0#U�gA�	�&}�%������߶
��+�9]�d��,J��oY����[�qk4�q���W�*�CO����*w�	���ȝ*�4BJ6���;5�]�_��;Ab��p�i��-��U�\^i7�̸���U�h�t��M։��䖱怕ن߰�N�xb(�𡝳~O�T����BwJ��2�.�(h|a� �: ��;dn��{D9`�i(���_���V`*���N���/c�He��S�
�jE<gn���<��p;-v{�
��UСj� ��N�㼮1��!"(�Q�h5eiѲfk��9@�CCeg2{����̂P��Ξ�;F���G������%w���y�6T�qbx��qX���HX���ϋ��Gwˢ�?��~�L�m����x("�v6)kvS3������q��ii���p0+oܾ���]|L�5�Wte����\���G���I��մA<�=�Y���[_�p;�T�\�í�����ɺN�I��W��� ̍| ��{�!,��=�а�F�U����=3O��R��0�ί��\�iƈC��F�K䇚��"c*�����0�*+Fx51�J=��&�0FSHճ�|c�C*r����Q�E���M&�'an͏��(+�1�w3<���I��l�Rಏ���)hR�[(�7o�����X�-(����
��?܉eBv�ӑ�PߞTB�ӻ����"���k�CX�Fw��I������/�^=IM���+$�(�xq���g���Z�4��ɋ4�ڊ̋A���~�U���N��Pŝ�.Y=$���I�Ne�V�#m�Pl��Z��;UyQ;?u�����a�x����5�LG=5:�o'q}3M�����\��b1 ��T�VcЮ!W��-��"��SЩ������x�t��PP�-���'����� K�Eap��i��inO�1OMkR������)`	�����o�'��ER���W�T�����������OC�P�J���� �aǎH/*���.,�4;�)���V�aag�DƉ���B:��<i�����Dq��"�>�U_�K��@3>����±l��n�#�G2�/���2���	K$d�r��s��|��,�W�(��i�9�3-E�WGcO{*���|�Z3W�óͩ�Y�sK�?)�.j}�Ͻ�R������g�H�ݣp�>�2���K�Y�nT���[u!'��x{�e�.�����bl���Y0ROl�w𚸰�n�Pd�o\H���RzFI�)�H�'��߄���Ĩi���ʗ��pzIb�z���8H��I�*o��nXg�V3�;�kQ't}՘��Ӄ��\U�*�:!&�+���ؿX���!�Xce/%�D�y�q�1�u����xE�_(�`خ�¤����0�Rk�y,��m��EO���a�\Bwq�b`�ݍ�ɹ����`�n� =7�*(D���)��s;�#�k�IM1��5���5Z��,F,��
$�w�r�}W�d�^,.��i*~Bk��Yߕ�e������Vd��仦>�f�R���R��3Z*���"?1p�b8�ME�zoUT!�1�ӟ�Α��JYn$��f��a�P����&lF���G������q���s�OV/qıf:raޞ� ���Z�_8��-�]����DI;�=!����o�'$5�_�|B���#+dC����ҥ��e^!���(��.z�R�k� ��!�O��!2��F���2���������l�V`_v¿j�~����FZ\����f�,�C{�ʜ��Y�]������*��ڑG��N|0��(�h�%u2(��S���-s��I	�eH��>$l�A��'�m=_���lAwa�@c��t(��9�*ۂ&o����IB���S<�<�<��l��o� 0�%�Zv��̪���B�`^5�	�/a�B����CЪ�cl֮�U�i�|@?�ʒ�ݫG�jNc�p�\���{��� �ϳ#����Wu}�݇�+IΨ*A��n�T!R$�_W�K�d:�ҋ;��"��Κyp��ߍQ�%-~pjZ=�2I��V��U���}3�>aY�m�l�v��Z���o��F��ь�u�	�.�x���ؐ�l2�P���?�HNM�ʴ�</K�P�NV�jx�9�:�2G�m��Ъ@�T�����D�(�Ec�!�eq��%I�j;�WeY��+l�ά�X_�з�.`a�s�Tu):*�5DѥÃ�C���ߏw!XcF�%[����I��� �
&X��e���ݤ[�wdj^��hG��.����e�:���ĆтIΜ���Bm�g��@��.f]��R)�C����4����"�\TY�YSQ@s�i�����v.��s�̏B��'��4�U�Xg�U���n��I`�A�_<W�>����(�+t���Ũ�2��JG��m�Ҭ?²�҄C�Y<��ki�z��x��9���-O6Y�>���k��z/(calA(��A!�U�J�a�n��=����o�����4x����;��I�j�ڪ�|c{�2�%H4�\4w�+�YD�++��%H��X8 ҽ��� ��'T�g���)S��Έ�>[iq�܉��9΢���5�]�=�C*�N�+���	X@���k�M�y��9~�C�k��G��ip-�o��B�7&<=}崣��JV!�A�8q���e-��o��0Z�b��cd"��*�`�*j֦2�}����������Q9|ZKݞ������Y�Ӻ��<��m���7��T�1�@q�.������-3V�4k����{n���.o�й:����qd75�`�'4ͳi�Eڑy�I����h������X/۬t�����,%���Qr�m��_ ���÷L��B�4x ����m�]�+�1
���XA�\�F�3�z@^9L�bM#f�e��n9=�v���� ���ߢ�8MGl��^�t�l#�	���l�#�kv�����&���J��[݃2�w?��C'�������	J���b�����|�'�РHΊ�������;��[V�Q�����/$���rJ��8�9�nM�C�{|ˣf�<��h��х	��7��"�&!�?�!\!�JP��s	t�C�~ڏ<��C7�V�L���Wb��*����~�� S%n��,�#�.�-��@���WV9	�7��T���Xx���x�#5dwq�%f���t����8 ���aV`;c64���C�	1'*Q��ᚒ��Q���.`���#jn�-������c�Qõ6���9���Z�#(�|8�+��}q3�1@{"~�RB�m%Y�LP>�c��Z{\�'��t�i( ��a�Sgd���:3HJW����o֘�0O0�=�u��$g�sS`}�{K��0�o�ر�Z�.Mʩ[�|�H�9$?cP#��%%��O��gT�QjLD%���s��;��ǫ��J@�#�����*��OY}K{�	�S��,F����������$;��+86�[6Iac `pE�2�b~v�u�1���%�����{ eS����L=� n!�0<�RID1�)��媅z�E
��۝+(�o��Y��s=�Gs�	͆��湧#�0�-��"��}ly���
��qLy�R�;�LC���P4G>S��O���M�d*K�kӊy�R�:g���D�NU�� �쾐ǣ�-`��A�R�7���X��w|+Gh3�҂�l1�GYc��3�������'�dSo����/z^�7k������ȠQ�Ss�Ch_��ݹH��]p�9�B��G8����g��\�OdRRk�F���p-��6?����Z�YL	UC�M� ������V��B�����ל��eŞH`���=ߞU�?h���В*q���D7˴L��o�ŎP��QBS��J��-y�\�Aȯ1�\MK0j�)�%�� 硥�/)�$!�g0��Tb+�!7)���X�be\xF�zس�z֟�#�\�q��8I�	�R������	7:oE11b�`�\{�V��K.�A�������P��޾��� �fd���}�ݣW�N� #��;�n6������0�aُ(1�(ˣhϼX��T�M��X�h0�?����k#8�O��3�W8�9N�%Ǒ:��F��-)�QF;7�D7�w��f��:���@M6n�7Zk#Q��3�O��+���u�AZ��4����-��&ҵ�fg���E"���cpvw���3�5όI�����չςn���촑TO����X�Y�\��x��K/�!�UG� �#A�JE�����	8�_�UЊ:��dK��HX�T]��!m��A(+ƈs��}�'�c�]J}[F5�S���^����nc[Q��_c�~4�*�G!�	���ُ��МV�ӵ,������9�L���3 ��d]�O^���\G����|�	��13-�#������Մ�!O�}@�=(�Q��PR EZ��@1<Y��d%����
�!�>�Cl�H6Q�Ka�`�"�8d�a�������o9)l�@L�k�m}v��_�w����ݵ��dV�����u���#6�[�L~c�t�Q�p&P��Y�\Q� !�)e�Q ��8�z��z��<!v�"(�#�pϚd�ɳwf\16P��i��U#���z�Ҩ#��`��e_S!`��ީZޅ��m����������P���%��L Yx�C�*����S�RH����a�}���|�$E��n����.g�e�0��Q!'&|Q #�Qs����'���Ո��48S��8u�z#�ty��71�H#�K�I�x�,��([]wa���{�θ��e�~��Z�5��&��O��;6�J���_��5A��M�����&;G��n�Z��7�3m�s�8�Y4�Dd:��yzr��΁3�BTMcwÊ&��qp���{a*�o�$%[��1��)=�WC���0���4�`���[�.���X/ݽ�C2�]l[>��nf��<�i3���aE3<���@j�s��&��	0m��/M=�)����$�1�� p����o?�'�9����H(G�>H��V�X4�VzVD�B�*�����3�r	��VE�P�*��z�#��@!E�N��m]���7i��i�N4�m�c؛��}���%x]V�H�Lvn{�}A���4&�ِ�5��afx�0� ����8n(����W�5��O��w>�[H��)\\B�iw��K'���IY(s�8[�:a��%}/pQ�ʩ�a�9Ț���$=�$f�8Pɕ�U�^g-����7T{"^=c]pR��CL�[P!�6�"#��FW�Ń���Xq2�3���&��Z�[��Ky����l�Ę\�������ʞ���N����gܽ����Q��Ht`�[�|��T�ǿf����� щ�{�L����[g�Y���7��c6�AGS O�k����P=�;�W�8N�9�&*:��/P�9a5O��S�0Ho%��x���s��Ж^_��;L2J�v�9t�W�M.e6d����t�� ��c��i��J@�BH�K��#Q�2�}y��ǱЂ��la��m�����]�ߑc��^�k�-�VQ�Z����a�`���+��-�p��u��񍔽v���g^j/Bx>V�0Τ��6�'����b;/�O�R>A@>�xm��ZΟ�M�*5G�Z�B����ӣMPU�؍1r���KC ���j����)h�YX\�7PR��n�8˭�u6���p�hw�8#V������5��TP	�k��:/ �����;���A��Oz�5���h�~ �F���G��d�)F!��U�)�a�l23��?�̗�n1�f��p2���XF���`ZJ�G/�R.�4��M�~�}��jh��ʧ�hr�M=��A�6���<r���P�B�֌�ݑT��d�*QUD��k5���M��l'��B��D�،޵o3n���%TSoc���)^��쀄�EE���|@`�2�]A����K�b[n*0���`L:1�H
^�qB����p閘��ٞ,u�|�t��|p8CH<��������J=(��l�ٕՙ��eq�pSX�d2��eqA�~K]պk����ǉ�RS��ڨ�4�'�8��������u8QY֎����c��(������I�"�uC�IM���q�Z��<�J�x�*�L�4�;N�60օOJ�H�/��lYk�N}�u AIy@�.	;��Z��٬��[p�\%.�Y�Ʀ[�z�Bh���o��L�Ϲ�r��x��g�*���U��b�R,�Y;ű�����{���~�ᐤH�,:�G���<ؤ'��*��ឞ`��E��VGs��M�ߠ����nU�R"�i~"8>^��;�1|uM!@w
��P;߰��#&"����2��3�a]8�rn�>G���%88�K���E��ӯ��	�_��!g4b�V���*]���H̑��P�e�<ϑn�r��C��R���#��ȫ��yD�@�Zd�b�ǿ���lbl(��K�ƾC���O���Z��:l-C~i���J1x���$B��~�kq��,��6�Y&�Un­���$�4����f�]̨�A�'�t�[7���Z+Z:��%���<����6*a�1����)>P�xdP���v�O�f��C�wk��R�#f_��hV�S���� �撎���#�G�9�Gga?�dqG��3��Y�	8=��}9�!s�IvZ��*�F�����-@�ͤ��l�e�f�b�3�J�'�����6$�,���#ۇ��7aH����h;G�����}<e���$W��aӻ'���Iy��"^���&�ά��ݡ�dPt�/1�(����m��ݯ<2�(�zZK5���+_Ե
@2Y����o(z��WEC��DJz׳�Ɓ����3�61�
4��4Z�$bu��m�8�
	���W0�_^��eE���@#z
��I�{�]�2�~���i�wR�Q�N�x����ƥ4��()�d��Z5��������-�\��i"�MO2��T��"،(�AsZ(�=M�l�x�)0Dx�S߹IPbLú�dw_�F=�9����5�*wi�JxI(�t������v�fEC�\��w����ȜC�c� ^l#	S9��L�5bo�3,��/��p�(��Pn,+��8SV����� �|�2��ߝԌO��=�"&^@Ȏ����`���r�`w����tw�FEeJt�G.$h�l�<v{t�A�%.��
#��^g	О�tݏ������}F͆�9��Rh��:�	���Ȗ�I���S|W>$w��%!6��C��f�y��$ +m�n`���%�͐��D�����
eb�.�����w"rg9�h���;q��5��^.BA��e_���T۩�:Lc����Q:����i� >D��$��	2$�k��"8D{#D������'�k_�!��D��A�FCB�.F��E�ҩ	�&�jJ��0��<d�:��rg�ԃ8W�-8�o){Ã~l�
JX���ՠ>��	��Ma�8\���yި\V���H/zX��_����m�Į5��R6���G�����x�7������4T�@��Lx�Q�b3�P++������2�;4�[�9� ��x��fг����Z��Y�F��b��/��.��I��>]�o�%��s0�_��&���ozi(���&��ݼ���ה6,�&I��|��O�ӯ8k�xs�X_r]�Q�A��� T8�TM�ހY ��]?R�o�'*��B>�m��9���ƍ{�I�$~'`������ȵ�'/�����411�I�B����_1�M� �s��œ�Hz܍�9�Ҏ�~��5��б�׷w�Q�!uC+�1�	��훮7��B����8���qz��a^Ćr�\��1�u��T����L�d�I�� G�C����n�S�>����-�/0(�\T����w-8"��DIY:o�n�t�����3l�'q!Z���vB�?�q�	�ԓ��>����	��Vg��6^3��+
�+�i�$Pﶓ�ۯ�L�<�Hk���8��O�(d�$y�}	���O��e����tH������� ����}�m��I���l>-%�a-���Eg=qv"�ض��H�>��%=d,朋[C�f�N�C���;���
F/!<��Ǵ�3/A�&VQ�yK�2m;�bHj�E�EK���3
p�Z���2��j1���z�!l�zl�AUj����Ș��`�:�X4&�<p�7}��� ��]�� |�k�Ĝ��mY+o+ѱ���S��.�I�>�&�3=9�����g���L���L����?�w$&bָ��t���@]�@^��6�Et]��U�����_�n&EU�� s�|��������1f[�R�&�(���~�Z˭+�d�D�/<�"�C�H9�*Fג��^����:��vm��w�C�Q����L��a��.E6.�U%�I���E�ً��
� �LH@��$�1�'crz�ˢ�<����ss[{b��� [�a����!K�L�����t�9A�k��B�"XI.U?����&��˰=x��|���2_�6a׵����믕��iB�(ű@�v�)/�S/f�V���O�0�|�
}�Tg���D]sC܍k|]La	�n���'�j��{��Р�������7���J��	:��O�J���P5�p�Q��î�Nt�<3�+��� 3�*�4���G����_w����^��}�F���{�n��KӞ,[
��2�s���K��k��	�GЌt�x�g��ۖg�u�v���Y;gd����������){��➘̖�,�V���{	����*���%&��)�ROQ�91�Ȏ�	+�T��
r�G?���m0@z7��$iO���Zd0>���4�8 f�|IS�6>����������s��
�s���OUu)��;4�� ��}
�{c~6(h������z�Bh(�px�-;�Bɤ�B�̍���N��}��i)�4�S�G������b7�d�T��pzS#�[G�Ʃj>�	�SgV}�c�V<z�\j�0����u-q�R�\+ҭ��DI��I@7
����[�ݚ����Ay��:w����SPV��P�p/a xLB�^/�R�}���+�{��p��2"�qg< �7X�w�-/bn�,��c�mM��(L�J�L%�
�VU�qk&y#�mY���;�l	e���K�{�,�� $Vb �Ѓ���8R.�Ϋ��A���Y՟n~V6�,���=[K	K�H�@+��u�9H���ک�����.:��<���hoq�p4��\udg��I����0�H0����%1�eߣOm�F�*�_�R�z0v�-�{�y�S�!ma�+��G"cZ ���f�b,S�R�+�t�P�������������6�k�*�����/!-I���<|/��=����&��"�>���7�V�e����5��_��kQc��� -~�yŋ��� %�Z6�'��eM�8�b�y�X	QI|/����`A�K\j\�f�\���K�]<�w�����A���s2�Y�^�祑&�����2R`�7�=���z��V8A=;	N��0;�^ԘG����X�Z�}<˧DK�#�e�UI�g�� #��t�k,��d��̰ğ�<ۉ
��4Nî,�q=Oj:�g�k6D�L���0{����nat
�:�����I/e틢��gx�����اmr$��C5*��8z��E�]�������[t$�؋��U�@f���'y�3�GOt2�I���.�@����I)q`���g}U�T�y�S:�x�]��yp�qc�.�zpL_�q��,�ݖo���#���"^}�񣹎��A���YNX�wjm���H�{�[�."p�2В���X'ؼ$�����Y���,�g���:ʭX�z���g����U���q���ig�_��Y�&_���Tq1��=/�+�$�{�'��^�?A�G;;��������^��Px��&(SOkmm�tU��}�ͺīv5	(2��x���XO�C� ��_A��M�2�����$�~$��DU����r_�y�W���e��1/�[s5�j����6[���W�"-����؝HY��y\Y׋�E�+�[ �C{A�
��z�@w+B��=��y�}��з�!�[��cs�%���p��t���}��c��c�,����<칅�S|s���n�>� ���X��3�$�Qr	��2�}��t�����a�Cs���fUo�q��3"���ϙ�Q�:����lH�`������EL�JjN�Q���
�|z�~{���;ŗ��V���#���a�:�O"2�8�.�a����gY�ƽ�^x�kn ���Nw�v�~���.�Z�j�P*����l�rd�U��L��XQ��/إ�^�f��(�oäY�JOmN�5��F�"���r��; X��ۡq�
6C���Ϳ�"�'MZ�k����r%mD����K_�(��޼O��XE�LB`V�N�9�)�Vij�^S�� ~Z������ʕ}�w�o��羿8�6%���*t�J�`+��ͬ��~�k;�|(�*���v���'�u�^�<��	�xJ�(S��c��»oF��6���o��J�Z��ɩa�xm)����C�K�œK(��D�s�����e������Q�B�\J��]t�[��B��ƣ	z$B�b�����cX�������Am9�J19�Ж�%���m�ʾGr�}��K��7G<���>v��>A�n�*�:n`V���zu���1f����l{��=a�k��L��<�z��d�[gi�饏A���q�Sc�'a���[}��`�k����5�F�R�/X�tl�YOp��#�n��:��Rz���
V���
��
��T%d��YM����1��i���><�1L��*�i]1G�!� ��.h�Jp�˦��ϖS�y_���/��Y��:�Ia�a��]��b�?�`�L���!�@P|�q��-=���� ��Ea�l��[>��mҙ�A�CQ�1oB}r�{C��W��X
�r?�|5�Y��yv�>p�sK�DH7�]�!8�I`E��i�5���%8�>��L�����H�I����0�+���r^
B�T��G�,�U5z���ml	f�Ew8�����<��7��߯��oy�V��M�˘3J��I"�)P 
�JM��Y�&.&��0�����#��$ʅ�&jm��Ђ<�I������3[�B� ����=o�s�X䪎�'^P1����_ ��'IW��6��D
 r4Y��11��QwHIά�	w�j�`�b���"k�$��8>|m`��:�K{I��M�7v$�b��G�h^��/_�LU���@K
��!�}��ܣ��:#�i1���&B��-��A��R�p^׻��Ta9��P-�m9Es:�A��t{�W�
��Q1�LX�zޜX*�gN���z-�κ�L����v"m�;9^п���$��춑ZGF!���[U�E�a~`	l����� �
���	7T;ü����dp�+ 9�&�����9�Z�8w��Uuh�	�����x���uB�a��� �L] H�1Lr��:"I�ՏW��):�-�>|dv�4"g;��3�
�����E�!I��ú ��H̯�$�Xv���2�T���M���+���yG�A��РW̨������ϩ�����IǞCk�[w{}!4dKp���EQmu�6M��g���'����e�f�'PS�'�{*�~��k����>C3ԘqJ�f���iEK+=��"t|��ɗ�)�\��xh�Z�k�C^�^^�R��nX�Svp�4~�!��NF��En�lNZ��lUvR�N��p��U����k[IWD,4�-�J*���]�zo ��qw�"����#���0�z�'�?�*���"1lr��̙�VLT���6���{�^~�6��u<�H�O"�-*�E:��AiT,Fp��v�8�?��{Nj��,aaJ����lnIy�^����t&��\���î��yRh�w�ϊW޻�@1��&����n�n5K����K����Ea�#(#=�`E[��[6���"�:b�9�nb�u�S��騿���kkи�8y�m��2�S��˧E�ϔ�*�?t�dNHr���T���(e�rH�vd�u�8�(�M�
 =JBUP�b�`�V�h����CZ�C���˔�vKU���&�ɛ0��En�:���/LV��E���x��n�Gbc��(7�R����T��-(l�o��&�ͼ��̻��Z��	���c���N>h���b�fۈDr�'��:�J�Q :�ꔚ���X�P��A����&sxk��}yW�}h���مV�uwDZhu����~y�����81^tt{cg~q
s~v]�ѱ1@j��V��<4����븯��`�U��8_ճ@�m��/@e����s3$"�Q&,�O�(�S�s�P@-�c}~���H�eF��|�$9��%�|��ś[��وij����9�Ŀ�C�����$t�% ܹ7�>_s�G&<��I5���x"����L�)r�0��V�x��[�e����/��������(��1�/��U�˭O#P9�D����JW��b���t�#NoA'��%}����� 98*�M��ќ�B��T�u��:������+��n���b�h��?5�@�� P�����̲�� J��	I�Mz�	�&2@aM�"PJ�B�@S�ҲDSL��*zR�����(>c��H�=
�{o����[ ��E� ��A�(r�%ҍO�ы�DJ ���W|U�ҪPI�����VF���r8��(��_��ۙN	 #pZ��Q���yY
��=-n�ހ�0��_��"���RJ���zh�3T+��K̝�-'Y��.���i�7�vx�	�
���� }���I~j������#�Uu�T���=��օ��ʻ�����!]�V�ҷ���&,����v#(5��Z�������9o�zۘQ꾡Rԍ�����쟤BB��Q��r[���.�)!��^����	�VySІ�K$��n@a4��!������B\�f�[hn�u�x�'�6e%���e��� �zh^=�L�w����.�Q�� 6��"W^���5�:�.��%T��a���vPq��9�g��O�)�(@5�H���Z݆Ug�v��Sd��@��Q��[?�}~��*4���������)�c�]ɱ��t�\E'�D��@d��-��.ך�R00;�4p��u1�!/LF=�59I�_���ރ�D�Z͂T�����Snҭ׶�t��g*��X�ť9�5aC+��G��1������~؁N��D��/>�l�1y d�@�'.��V����)9��|Y���p���%H���GN.�nV�,�	�i�W&+*��K�a�p`����r.��It�*K����9�yGTlԃp��r@9w�G��<тROy�:B-$i*�8�F<x�>/���A՘cҒ6���|� 	0���91��"��)+N�-V�e�	���J,5m�/��<�������t�Ͱl>��z�w"��a��:���&v�����7�3{�L&�<��:FB��d��bs��7�{NCН�g��r;\����?��X�%s�t��_��ch��c~�J(�X0���F�X��!H"�'�����u���:#�o&� � �3%���.҈���`�p�Yz �uϹ����fj�Qi�b1�-R�m�Y��gh�w�N��\�r�����`����/�wEAl�~1w����Yޢ�E7�P<mY�/������
�(L*�̻���ҹD��5���cu�P�weGU�&J�[{����g���c��.�5]�u�E=(\�STه��"�{a`�ize3Q�?5�Qq�^'�B���d�7��A	��^�<C!��f)�9ɞ��@u���2{Gb���\��YT���Q��8�}��w�7�&\����"MdOl���C7Kyh�2�y��b������13`�,UF�"�N�(�t;1ƅq������I����j�D���hj"��C�!�yQ/Hm��Lv������K��3t�т0�Ka���m���1TP��98p��u���,%�������IS�����YB�VF	X��ag�: ��g���9�O���rUw�*��,�F��e%\l���ZD`9R�Zi�&�/��XmBMX��&j;䵧�K*�Cf����H�l���L��&��)5�\j��Z	��95��H�M�b{���B���#�����Y�0cO0��y�s��\�T/�a�Q�"��B%��e�F�� >��vyq��X@�z�]q�)���0JBXy]��qD2?��TH��ϼ��kPY˺xh�z���y"���IR�يij�E��Q�����P���ņy�}]���z�cۃW@,�&D9�zz��Q$>�f�d�`\�(����u� Gꚾ̼>ߐ8�M�8x'�"P�ɕ����c��f �!wr��-��/�-;�'��R��I߸S�Yk�ZQ-S_���pV"��R�Ȯ5��(����J�i!ìY!]�%>7O�@N	�m��w#�q����D�8q��وZERa�����Lv6QVc'A6�]�<	��p}H����~�H��r�������C�K��<5�N�eb��az6��E>I�t�*z*����3���6�].3����4�RvQ�Y���B���1o�7��׻��dΎM a�R�L�Z�i���r�		Տ���71��Bh��?��E2˲8�m`s������lJ5��,)���)�zV-�~1ڠc���D�\q�^�*�e� �c_n|`����W�m�b�u K����Q��xWY���9^٧�������Ί=��6����ǓAz����պ���YeB?�(�!�2:�l8���X�G�iu�����y�>�z�1�Ĺ1?ȶqA?�Ȓ�?�\�+O���?�䋸n܋D����΋ѴH�Ѷ��O4�bs&4s͆9I��-0�,������&]���j�|�0 ���v[#(d����$�R�tL��6�5e�&e�d�u�U9�5u#��w�h����4'T_qAv�mQY�]��\Y��CF��z�Ɇ��4��C�$aL�[�[{!��i�	�C�m��9Rq�Y-ӠoOz �ɠ+�|���q�����Aƹ:� ��A�Ӭ�_0KO���XN��š`o�t�b���L�/aHj�11�	��w��SeD[������惲ř#7����m�s��$($�����a����ݦ���}����z��y!%�R��)Sd#ws�'���l�֡�i�\��c�D
N���� K� �{U�`����Y� "��¿J��u(J����iԝ�~ ���(���ã�a1�1!H��������w�2n�3,Md���7�S�v�F�3j]�J��<�6�G<��D� �	~.{��N���ط�Vk
�H3��ޚ�RT7��Oh�Il�,;�v�G�j��� P�,U�պ��{٫d[(4A,�C/�>�{[m;l�xj�ׇ�c�/� ҾM�	�G2���\��?�!/�'@W�P����(C_��z�yvo��ĕU��=��͖B��2Wq��������`>̓D��֟�X� �E�;�g&��)�&�n�:�f��U�lq�y� M̸��趓�.���qR���X�H.{<E
�s�@��A���oQP4$�'gȽ��0�B^X�U^ڂt+�	F�u!Pَ��R������~k=�>���4�7k�C1��)��r�ǆs3\PMy��*����֙wJ@OnM���2�+�����M�ǭٻ{�^�d~��s~��ݚ^���ny���_������V|���@�]�����'�L��!wq(KT}��
���F�]]�_�0��#��C��
�E���ygX�z�{���ĸ�����O�SЊ�X�<QDӑ#P�~bq$�������)�>��^*)Md犷Զ4�r���6��	�V��U�07;D���p���������~�K|��x�n��D�4����|8��IF��G�Hܗ1��Y<2�G���vfk�7N�v����1*!z[��Y��<Y2�=�͒#�#��S{�v���w�lB�N�+ң�SkGK�c���̚j�%R��&B���G8Jv�j|�~��Qо�	�3I�Uu(,O�$�/�8�c(��"�g=1"������ar*/~XJ87�ɇ)Q��]A�s�{'-��*�G���6\�f��F9|�X��w�zOB�K%ާ�����y�g������R�T�r� ��y]������IX0g�m@nyT�/�:+k�R�/�7�u�i�މ�IHD1��<��z�,d�0>��T︵����T��9OFe�p����n��6�j	vI[*����^p�fq��&��rF��h�	
iB�Gq���/��Κ�5�DA"�@���鰈���\�0!`}-jr��i%���4����wh�F���:g�oM�enq���Z˙��b�T�lE,��k{�EoY�"�7 4&�ψ�i�`jQ�p�t�����\��i�TX@S-�X|�j"�^`�p���7��B8�H���M�Z�o�z46&�鑅��<8�@��"����/�ʝ�2ܥ���<oj�i��]yt%"3ӟ�� ���m���/���f�"g��R9��XѦ_*=27	e0} :d �<lwI�A�a;;Q;��5C�L��E�2v�<����NÜ*�7;IQm	a˥�v��ů Ս=��~l1_�$��Α�S y$5;�sFُ�p�O�R�����[x�%��/}~{�H���B��S�l��ޫ�OmΨn�,�.���~��rE�gu� A+c[hA��,
�f_ŵ^"�O^^�0hڄ��#{P�1unܓ �h�J)��F
N�y�2;	\+��x|[Tvq��
!�e�a�ՙ���쑕g����gp�����(�����H^��ʍ�1�C8AI���������7m7��W"6��Šq���߃��[F�*쎡a���W��w[`z9ϟO��3,�1�����럌y�l|���y��| ��/jP���y�F�
X7S�d���#Z�>�Y�����У�$�t*Q���C{O]�*�ŀ�S���ڂ6_ݒQ6���v	�
'�`�Ƙ�S]���+~��1��o��TAH�������ʅ>�a�e\z��d��}'��vQ'�g�kl\����}Ӧ0��H�����c4�Oa(�ɚ'�{�%<��O`!�J�R;-�9^t���?!���k�����\?�}|��3�{ ���b���k�Pji��A-�l�v��_���P������XZ�:ie`��zS��|��4I��*}�B=�r3E���=D7��h_���P_J�ߙ|�A�u�T=�f9�D��B�| n���dv�G ��� 30&�}՚\��tM���D��IG��#�T¹/ܴ)��΄��g��Q����;[_^ۙd��f���H��J+�Q-���U��	&)X�*�F�G�5/��[]X�Ώ��00���[�!��4W9��ƿN�kh�y������ܭ_�&��ߒ����H��£+�XWQ�ѩ1�=7�	�r}:�9� r��,/�60{7�oq0�oh��#�M;}4`c��s/��"�ko�~;�:��cX���[����J �e����̭�0uل��]E �M2q����D���r�6����/�b��̐c�P!4xŊ�|n���*��=���r�Ȥ�օP{3_ZZ:�o�>�<�S��7�V�u���5�T��s��`7��Y��%Hl����T_��tQ�3�+�A�sٓ���Q�=���]q�ps�
m�
w���� RN�V'�&^L=ֈ s�l8+����\���E�8=|B��r�ͩ��H���i�$�$���"� %쩫N��@Ќ%�0�e�u �G��x�_��)	�p�]sμ!�	m3Ś�A��jiz�aB>,�\�5���E�^�L�A�{]V;��j���'ʉS�t��.""��>�J cD�x�B���D��
�<B����[�`U:q:L�P��u�6sTYnƔ�V�|F�H<x�>��eXGI@�Շ
/mf&Q�����R��ۇ�G�3���蹇����Y����A`�����ڏo~����χ�ҙ�w���8��n���w��^H�w�e�]k��Hü}iШ+A7/j*wc���}�%����&��)�����ӟ�uI�զ�Ue���9��y{���Xim��&��c�HQ.�3M��,)��F���<�+�X�������iB��#�S�Ei`n��UEZ��T�L�7����ҳU�nIY^X��~���m��x�ʹkP�����FiY�4%q�ٻq���B�ć�Zqw����́��;��A��k�]��j��(.�:�)�Ȣ�&ܝ�ڙ�&!�w��P�IE[�B&�KE��u�Ȯ����Q�$z��g��W[�~�����(S�3�wC������J��q	�fE2;k�w>;��GvP�ԟ�u��/��W�̸F��tq�\�A=9�e���P�ϋ��!���Bf�V�M5SV�x�nWSM�;�B�yo�5��4*��%�H�)Ǧ4� 5��D6���/�ѿ7G���1mˇe�0"���׬+C��1�md�Y�T��"�C������Zx~z0	܄���)&ڲ	�+0	z����}��]�o�A��=/�e�Y��{M6r��c2�t\����AwZu�V��"�Z��Dv��e�<5S�,��s=��S����1��k��z�?��G��PsÁ�R��YW�8.R���>A\�.I�_g'8$`��8Q�U�"�O����/_vF���'��S�c2x���?ǒ�b��'�J�[]������H��}r�Z|����a�0�u����݀}���#�mخ�5�&��w�=���L�{��x>�=ɸa����6C� �y�	��CxNX8(B�Uv)���q6bn�9�.]�r�O�/��C�KU�N`-<{Y�@�2Ԥ�+�E����lS�y�~�4�k ����fIv>[9A���ݖk̪<�P ���w�y������y��;F͛��`�)t�����|\���0���e_f {2Ij�PL�\�0�TY��|�ױ>.M?��80����b�Q�(�*$.�=D����<�.���G�B�v�~=��!��[�ɵM�����$X�]����G�jMWU�5�-7�}��nt/��Rl��noԼ�wo���E�Y�'$rk�や��������N�xغGRs/1ymݮ\_-˟JE�p<�ZO�M�`�-���ēX��=(�ʮA����C Xg�O&����J����s�
��a���H�Lp�z� g�P�_���mj�����M+�h��"�'�����$/��>��g��rU�	�����rz�&�DM����r]��]�@�Yw�Ƹ�(g�_�g^ӕ����s0�#�Ӆ�춤w���)�lg�����evey!���9�h����C��r�|������k�@V�_
}�nEF|����%g���%M#�ʋ�uM'v��Ũ;G4�%j�O98N?�]1�&�
؜yأ�j�l�(�aO��B��o{��4�r�PC?i���3���fp����?���f
'�W�J��ͼ�\T�x�#6~1���@Ph#j~*��լI���Ę�U��Y����/˽�O)]�Kn�C�� _��r|�.)�(	VI����<s�P.��*0��4�-옋�]}I�Z	��pZ5�����	���������)�Z������
q�n����q���n�~�W`_#H--k��b)���zϑ�mL��Ɩ;cU\�77�,���-$�?O|��-��S
k���2}!3/נ��쵾ߌ��X2x�q�C�r#���Ho������R���,��.ϼU�_hv�Ad$����Ma���Zpf!-,)�Q���0:Ɓ���~")H��$˟Dv�H����wz�p}��M����Uo�f�����5�syߞ��3�yz��&	J�̺�Z���SİZˠ=�Mh�D������S~�(�D$W���Y/�9 �|]���b��֪��LTB�l᧼�L��Tƹ�zu3��dB��	&ܗK�0�ժ�c�Y2����D��1V�P�0�ig=�*���XWR'�X�t�Y��*qÀ����Ga$pt���c˔��X�|dn� �o5�W����]}&�?m�y�-�����C��J����oT�V#�D.wu���7�_d	@�_�l���So�([h�U����<MF}>�h����q@�dx��.��p���q�1q��*gh�+�)\�O�f��m�m��/��50���`��oT,��*�?,���ߦ�"�w�0<z.�d�@�\�M����5\�B��N�g�i�K�k5�}�a/=p7�j=��^�H���rl��s�Ӟ��J>���~����N4s#V����]�p���"1P��֎ά�>
.<��ʫ�̝��#���*�Pb����T�0Dy�߻h�����\A橆�K�l)���Yr��X��51F8@)�j�X�Y��W_:��0���LL�<�B_8ޱ���П����097�N0~eb��3����9��L�Z(?習p"��p���F�uOo�y �e���WY�v"">^N���w�������7ۻ��ۆ ��f΁����SM�^�(-�(�t�4�W�Bh+��m~�k�4�L�Ɣxs�<��Y�fM��C$��*'�{i&;x��w��6����]���o��x
:7��(����ݍ	�M6EU�A�<N�ZX���(��º�\e
_e)�3����N��)\�/�ꦧ=��c9=&�_	تZ��n�Y��D��-=�a�5�D��)0���0�3~�2�a_�_r� z�=Y��L���^�I��~�K#Aal����I	ǿԯp�o��e��w/�~�.L`	�(��)��Zg)����E@!��/s�Y$s���1�VR���e_�O�)5����%lo)W\�r��k��n&yLI�,��،i����G�N�[0M���uR�ۃ�*S)��N�:ice@�ϙ}y2��(}�Tk����p:gV��Rڂ���AD������8iMH�Ui�U�m�I���D�X�߬i%B��P�Y���n�ww��^Xp>s��gا"�̨O�\�lk��@;YK[A,�ץ��F���Im�t���f��[����!����nEB���$,�#��#�q�lKs$�C��6x�yM5�	-�����~�0'�a�ie���(��!�TWp)9���|��	�`t��(/Q�5D]��B]�y�6ٖ���?e�P����y�����,z� �Z��2LC�u�u�ԣ�eئ�JF=e�@D���9s�pZ4�N'�x�)��з�7?gw�D>
h�-�Ŧ���8�.�?sW⓺�O�m�r���F�G������F�u&���y��9^�xm�r�P�A�iۻ��8�=�_f� ԛ����m�PdyH��>猳
.�&o��>^`�0!m�g1�'$ؔ�|���Xwm��u�b����\/>^@I܍;�����o&v\%3'����\*Ԡ/0�󤊖x7vJ>5��(�w]�(��F����LŞO��X|Oq[!�ګ�/jLQ,��e�p��K�]1aݥ�XC��yN[�+��O�Q�iװ4�0���탼�5	���16��$Q,O;��M�����,J~�X��}��c�x�����a;��j')3��R��#	�������LR�yG��g�K��y{^bS����~����k��#��\2ߜ2�N��!�u"��N�9U}:	� ��IT��N��	c�glx_��nX;m�5�C�	d�_�!e�:D���i	{�Ā��_�:����٣
�FHn}�����&L���fr�q |��.~+��=ӧ�/�:>u1�}�/E���o���=�LiWH�p<ee>���_� �V�D�5�c=���brx>a"�z��Oh�~1���G���R���^G"��0���̇t�c��wYg\6H *���DЫ��f]��Hp��fLs���3����;R�:�RQC-���t�q�T�s�����{f%��*&��f�0˩�D����'�t%� JAڣ�F�U������s:V���)�E�i��p�R�!�y�g�+����9���/�d�f`�_ը}&kT��"Z ��C9k�*4P'#�w�Oɂ7�����e����;UFH��������:�6_f3ZN����9w%H2���bs<G�h��YɶnO��-�sȓ�}���:�BX #���Hq#w�ǞV��M�|Q�B���3<�޶�O:��%�6�k�?[k����d99�s�&���3FC��(0�t����̯
��&?���KŇ�s����B��Q��^ M��3���;��[�z�}�΁{��ؙ�b3d��}Sһ��������ו�����Ec{��⸆���`���I���`#�м�N7ޟ�+��@:Y5��sΆF����֢q�hқ21��WҞ�i��hJ:'�,jx1�L��<��b���	@�n�6��/N'0 �Ȱ�����bk�����b5Ef�9(� ���ד�2TO'{�cN|:�#|��c<�5�AX����}��G���<�r�}�-����9C�6���8qރu ���r����J�!�j��Z(]!�{� �F���&\�e��J0�ޙ;��b����P6 �ϝ[����5������O&-J֒�"�؄��B���N��w����k��.1����,xfױ*������`��(`ö��\^	`�}J;O�25
�N�S8��d����߉X�t��'D��B�	$���)R	~Ƙ�AovcŪ�Hi�u1Ww��K5�{��j{�S��P��X��c!p�;�9�J�.��h���Ѻ�" 1���Q��գmW��u�A�E����Э��*⎠{���Ϙ�W3Aݦ�Y���1��L)Q'��	٩�:Kw��0��oz� �������X���e�?�x��W,��x���Ӫ�+����D�y��P��KoR��`Z�o1����A�B�C�H���V�H�~T��j]f��H^d�R�F�k� �f��γC���7g��)�- |�aq*ݻ3�Pi�q���mzm��$}L�'���Qf�x>�ge��O�t�>�v.���ucơ��.�����6Gd^�Pif[ ��H��lM�wb\f�V��Uz����-.��[M�m���ٞ�t:���`|}�E�6�/Q�^0~�s2u���u`�U�m�h�Z�=b���M��8�c�ҵ�P�2��MJn"O�:�c.ˇ�j/Sf7�D� 8�	���Y&�8�Fk����&M���?l�w�a��[��2g�p�]۬e���Kv˱�@��]��г�5��V��@J~��r�	�e��zJ�ĵ��;���+�0�ݘ�0&��D�&u_+A#��L+�<��PY�>���O��w�о�?�8e.CST���kG�����q��/8�ܤ�}H�x� �u0?sV$���B����\���ɲM,DGq��v��|h�h.���N>^_��p��Rk���2bU#���*x�e?�}��ʡӑD�bl�;�`��<$*��]N�!�eY �˨}���覮���a��y�%W��_�?i� 2S��dU]:>�f���;�h8�R�`,��qy=�Dd� R�,t<Fş��Փ.*������
g�_�`��e�!��ѸO����-�[ҳ�]�[�/qￗ2�4�s����@�-��V\e���"+�?%������ŌCA�s�3�GvDlb�!������*%�#��>/2�/e�R���W&*�Y��;��M0�$���*p����)V�ꮼjd�RREQVvc+۟�n��$.Tih��7q�N&%`��ۣ<y�Z�%v�;�Ȓ��.�J�TQ�-�aO�U�Xd����ҁ����z�*3��s����E&�g��Tb������fs��p��͊+	嚻��ܻ�+�+�#�7(��yc�R4��k��G/�if�	��~��N���C1�#)�OR$K�E�">'z*��d[//�~S�)}y��*d�wA~%�V�r��-l6Kx�5�DS��0�ͽ��6��{�;5�_�]�܂��������NJ<W߱�ά���4�fh]P��ÓU2´�=�D� ��@*K$����j��f�ʫ��j%%�(.-݇?r��!N��ギ�P��q���:�Lx���ɔ@K�C �+l���|�l��E:P�>�~Ovo;�� 6�>:�(���P"��ǥ,Rv�!^h�J@�Ң����3�%�Ė�k�lj����\�������i�1�(���=�5��pI�w�MO�K�K*��uOܥ�n�O �/80��f+kH�K����W�o�<3�OS�Q�9�qs�?2T��*��A���S��%�w��Kk�F^)�$���j�>	�@
G�CY`E��G���-EW8͌2��cXD������!٪%�dG�s#�$�k�Ra�_�Q)D���YY���@�����7 �s��E��G�ni��/��K���7�sE��kA���,P��Yi���Ā�������P�ר$O���J�wM��)�p�U^{oI�D����S=����:��,v v���e9���[��ECK��k��@���'	@MV�Z������n�������w��}�,�O�5��[<�g��L&:�<�ܹ=�g>w^
�!�c�M%��wbL�q���5�I#˒T�ڇ���|?��9B�R&~�N�@Y+��E���/m�2����륄�=<-mD{�CX�;��E����� �K���+w��,�ڎ8��R��	���	�	r�ӻ~�~~$Q.�C���N.��E�;K���z����}�1>w�Z��:���w�4N�
 �ǋ�@sHlL+ഘR"Z
���"bJ�1fJ�#�`��Xb�*C��[�R�@�i�/�B�ߘAk�p9]Ƙ�~�v�	���/�u�0^[�	��ugWw6
yz����
]:����$Ɛ85��<w)g,�mN�
�\Q�x��?b(l��ǉ.sA�Z"`H�ˉ������Sҟ��H��x�	t"�ĩX�j��m�X�Vwj����"lU�d[�YWd7�oL�9(�igg=�b�V���A��ZeymV�R?��F�ZRO�c<Sf�©o����܈��= �]</Z���8�Y~��o������T ����8�u����ݞ������Gnr��ny!:�-��u38��_����sQ��n�>�5w�t��hu���ƙ2j �L�4 �8��kp%�;��n���y��PN�kfٮ�d2�YRt�Z��x�S�6U�F]��(�D���,`ɞ�(Sœ�����-y�0f̵��H�0lj#���ć��_�{���L'��2�׎)�7�x#��@wkWP���@�_�K�Y��5q;�H�m,rd�TE�fnڡ�N-L[�&�@V������B�fqMҏ	��}i1����R����6� �:����Ȥ�Ch*1$<Md�"	�q󬵙1S���+�Y_Gh������H�w=�hS�t�M�b�N9�'O~�V�Ċ<_d�H+�Q��G3����Y�m�U�Qs'N�'�*��|\����	5Ȭ e�eC���5�����U���!�-U���8>X��o���Z��]G�J�X����dWn���u:����w�8V�����qD��8&_ڍ6Z�`|ڑn�+��߶d��xn>A�8$���bqs�ձ ~��t��60����6|��a���o���R��#sB'?J��o]7Y��5�Q�|��x��܏<H����k�J���~{t��j�9H��L54���tQ�?&�	`{���rS���K,�OK�J�-!�.��p�z�Ϫ�ݠ`��fzϋ����J뢚y�C��۳�-�4�&ߦ�i��u�?���qV
9���:�O���G�r�� ��G7�a�.&�hZ�iX�T�;��s7Eb��6>��mNH����t_���n�����ٚ��~�$�N�ۓRf��Yh綆���`�Z�V���Fj�B���*�m"�{
�\Q�4�����/�0U���*��]0=�;'�M�@�qGk_�vo �]�I3I�y�1��
z?�+����:gtg�����8qHV�b`77O�
h��;��a$,������������=��% ���`�x���tCP���4 C_a���=��W��*��'	K���= )�v<4��c�8�f1%��XwBU�B4\�'�r��+	��y�_�s�6<��^��Lٗ%�5���A�:S�z�J �p��K�6�o�����z����$=6�����M������Q�>�4���Uт_͌�Ӑ��������ah���r1�J��L.����64L��f̘��gJ��8�Fy/ˋ�1J�����M�y��q���� &�y�8��M�j�%�ʅ�
ƍ"����|��E)8@SL��D-sx�f4t<a���:�N�I;���,��v�泶�E�^_ɻ_��kӂ���U��.��5�b��"�uQ B���xL>��&l{(tg^�)��C!h���o'�m������M�t��aC����den�'L�]��:O~�����)���ʴv�|��$�`�+w�t�@�C�1:�6!��xtd�2�tr��,-���8����_�$�܄ho�C_��:���V��x�����Lo�L���3�|*(aJ�)�?�e�.�Rf<4ْ�A]���Z>�w�����������Ɉ�qo�=dw��.����FYi�"C��s�J��٤5d�dR�.#wp�!:����@}܍;�*E�#O?R�M?P�-X��	Uxm�H5��%�~ �4�-C�$8�HAj�s��N�x\/�d���	�Ag�bD�o/�ym:<��K�MK��.vpmc�.5TwE]���+Y� A��ʳ��o�e�|�M��2�9��Iq1�'���u���6&`|j����f��;R���ƞd􊬤�V�B���������}�.H�3��Y��?ǆ��M���sȺw��ǧ^��C��tpɪ��.k��o�R�*��%�<�{�!�4�H嬊֎ٻ?�����??�W�{�8Z��~dq�2w-�g�o�^gP��
ɫ����$ь��=Ǒ@��}.��xtcʊ�J.�=>L��cM�vq�y}AWr�{��,�����F���@��jѰ��@Oқ)exY���$�v��UÒ����^7�[|�V�����+�ρ���>xv��v�>�z?T�9�R77C<�(��JܞK|�_C���M��_H?�:f�d:w���b�8�w�C��{~�?@&�yW)Ъ������$=Z�B��GmGi����8-|V�>O��ͭk�$�К~�8����j������
) {=ZjV�bY�s�ucԋ5���Ea]c<�𻀣�k?�������W��#7�o�/5�@h����I�c����	_��zu/S�0�Ƽ����3�R�R�z~�g7I��AZbQ�֫�<���ᢐ�%uם�
Ͽ��Ȳ�+-�)����&�A��؄c�}D��4����E���ui��d(u�9n�p��iԄ�B9op�^�����~�J:��ps�WB�;⎔r�f<�id.&d�A�%��Y0m-ʲYqػ����|e"���-�h=���dSS#�l>썟̑Qt�4�h�*PO7��b�a�6dI�;ߛ Q�|� �=��w�%8Z"	��29�Z�w;��n���3�����@�z=9<q �ٛ��(��K����}Ǟ�D7�}�|�<����d��֟�&wW�����g޶U9��N�{BZ��=xX��D S!:��ΐ�yp�/�ˬ��1H�9\eu���(�q.���Q����1�N�7&y��VR�L���0j��r�_�O7h�,�:������ot?�dm�L�iWA�ԃ9Ѻr'�����'/'����E޳��^���=A@��o���w�\������w���W�Ү���'(ƶ5�(C��Ġ&���W�k]�ſ�[�k]@��0��5
>:!�"Rn�b_����kQ%�T��O��!V��]d�
�4󎼙ی��;Eg�ǿ�&Ix�brgt�5a ���d
l+�3d��z�|�b��\�1���e�Ĥب�%����f4E���E��y�^6"U�.h���i�r�-G��������gD�,M��9#/��;���!$��9k������QPiz�W)�ϒ��4*���]�"9R8D+Xi,�0ro^T"z��Q{�O�̲W��_$�G�J���г���
ݨ+���<��Y�;e�t3Jٝ��ڙ_�P}l>A!���'�/�2�b��ہU.5/F�yR�����(�9����-��A-�C͆�"����B��@����JE�jpuS|-�8�J�@)K!I_cG���PĲC��h�?��_�c&e0�T�,l���q�d��4\����K�8����o𻢺,�Wz��L9�p�#p�����ӣ@z�SWM�#Ӭb9�M��5���V�
JP���Ch�Aq�F����[)[.��i�� ϡ�'�X�#�YB�*�$�3�~@2�ǰ�c�S��U����6���&5B���,Ҵ�L$7��¨�:3H�+6���AW*��X��9�L��r2�Y�F�7��c�_�$��wsԼJ�㳷L��Ar<�<IۑzPyn�	��tD4ц�L�	�V߻�@^E`�>;[.��k�u>�}��0*?F^@�%A����2��p�lab�ZY��$�{c2�W�sl�:X��ݯO͍�$e�h��e#6ŧ�D�'m84��^Aw��x�(Z-���Ak��H:_?=�����Ŕ@G艿�UաW��Ӎ<j�-�Q1�ԟ[�:!R����h�mp�Z��6"x�����,��P)�/��L� ��˶�i
���+�w��̈́	p�a�����z�"�m��m��E9��rZP��?S�T]�6��_�1{��fm���nz�l9�t]�?J!��� �>��������b�>�tf`[9�DTďϛ�d�.�tǾH0�<\hs�7��X|�y�6�d})�V��@���B�ݞ�p`��n5��E������B��+{�.��b0u��O�8E/N5�5\5����s���Yn�D2�\PJ��5��:�D)�p�h!��!wT͚I�v*@�7K�ǆ�S�T�t��ɶ)��5q� �����K5��yQ_lS��Z吱<cP��W��;/9�n^��ɾY�ݗ�Cvx�U
�e��w�߳b�5��։/5;Iu	�h8Ѵ� L.�Iz���Aah���~bS�ڦ�¥uc!ɚ2G>�,����P�
�;?��v�0f~�#�'��^��{�b��Q���6~���db�wR곈/vQ��nd�d�]+�[d��/����f���_,
.��dx����410�3�
����_�?��^��>1���y�f&e�������\
!�Q�Ĕ��F?o�.P�D1��"?�JR��������\]֢��������:?���s^	�N�ںz4�,l;N��Q��ل�Q)y���Fe�!O�hݧ�Q#����o�X	��#����耈�]c�����:"mf���) 6X>��dg��&��OJ���r�}X	�����+������?�l�����6ʫ��qUUr+�t\bZk�̩QW��\�5�Q���g@P�:�a��J��{���� �8@����饅V=m?
?[�	I&��I�i�<_	p-�<>(���� �6�wLU�n��~?��M���hQ˄� ��;���������9�E�4l�X���%���t��I:/Z h�%澜ZvsG�#�Hҏ`���Sg�0��'�ڲ9�y��=���#�7��8vv�s�܊�����zZ���4�Ȃ�D}i��y��W}�:�|�}T�|�����S�Yj����,�S셆񵦡�⚵�]<� %�Iҧ#���}O� {�G�"�}�Vcľ�c�.���1s"��?;���(�z��;e4VT���9q�9��@�=���
���<�`fJ6����n���j$�ʜ�4wD�� ��\�e�I�5=���#�v+��d�]m�
d+�]�)� ���ߔ��枧u).��;��|!d�DK��R�b޸!��)�K:��+�{���6�a�s��ζ����i͓o�OIU�L��%P=t� �;k�T�˒���,l8�dlh���Gt.��>��A�G��,��e���ۈjr	&Mʤ�+�WYc:~Ԟ�-s�h�G$p2;��$�}s	��9��g�4�4(e4j�1U=�T~>:w���p:AĹ"�g��ӥ���Y��ţ�TY�~x�9 �����䁁��ɼ[��0�4�@# ��Ʉ���d�/�ܘLi����D���Mo����:dܜ�xtsì���j,-n�%�&���߽��	�ȏ��jAO.f�d��ԇ��ǲؐ<y��M�3xk$9
���4*,B����:Y_�R���z��\���R�jZ�2b�Yz���ΐ�[yg�W -KPF����F)��6%
U�Ǽ׬8(�2�-�����	����!�wg7;[�V��[I:~���P6��+OY��'���X�n�a�ط2Ą���)����S��Gdn���ll+����-5�Q�O
q|�GO�?0w:!M����UM��%�;�� l��FkY���)B �aD�b=w���F��R6�TR�}��a�z�r�Vf7S��$�Z���9�Y_�H�B\D1�;l��w��ox�}+`z��R��/��n��,B�4���ծ�y.]�}	[��猓�&V��q��uJ���h��kTy2G�%��a�^��mUoL�H��:0N/Wl:X�wX��(�n��s�����~��q=^�;�	���s%pҏsV�ŗ�z�����Ga�3�p	z�T�vqǛUq:k
�lf�~��|P��r� �{&7a�;UO������#���z��F�؄��%�/�&C�1�ˮ4��c�C�zs��S�J�+�/�ie��_a�ʄ�٣D��3wBﴫ�
9M�:t���j��~�)��OB2�93��d��M�YǤe���׽��Qx�c)ݦ��W*�_�G/����� 5g䜕=ECR3������o�!ח<r�p�v_12,�tKfߩr�Ό���uCS�b%A�d�"@�VZ�9���N쥔���6riL��ϳs{�P��]�߅9'�l�X4��{Tpvr�pƥM�
BF�0�9:y��'	qI��K���>�05�c�QC���h���,E;3�ڛX�Ѓ��
����?�?���ߧp�" WǏ#O�ቡs���	��fvn�U����?�|��I�о/FrJ�VM�^��U����^[��<����~�Rawxrh�c��uOrZ7�O)����I%�rG��gއ�Q�­W��j���k=���V�%��ז��ُ��?�bR�Q�R��-��*w�.�ر�[�k��'���*��9-=ӗ�1��29&�qD���n+��S���a�m����@��_uܡU��[W��қ��;�{}�e��O�f�,&��W�J/�Fb��s�g�@1����v�OP<z%2C�/�g}�cO�"�ʓ���l���.v�b38Cw7��%Έr!�M���������lQ�d�d&6ʒT��X��ಊ�a=j��bI"=;�=7�T:�\�]X�Soh@�0|���-��hK�l?�:�����ElÎ}D��xP�Q���������Vq�\p��k�J	ux��]_�sC3{?<�:�������n�h<�}�$�}����hI��%|q�)�E���߽H!�r��N�䣅����/�s���u&ȩ0u:����@@K�/���m���E|�z[�ǈ�=;��V�K��K�NX���M��g$z�:���0Ox)+�U�P_ߟ�F��灺<cK���B@dG�"��;J��F����g6���jX$�az\^�t2n���dǪ?>Ź��1�
�Z��*��ҩs������8��n��퓠$뾛�vQ��{]ƒ{����oBGX���J�	�u����z��?��S���LN|f~Ó�!P���z]Vf=��_o��ᮍe���A��M�C�a����4�j�1Zn�`G�'1�����_Ȉ��V���iE߃��	��s�M�\0.@O �l>A6|�3��a,x��N4O9�:�0��P�7bvu@1f�9d��әۑi�+j���!B�YI~ ��U�F]���X�)�B|�s���_Ū�/��A-K�l�0���d���+��B��x3���Y{�n�O���a����'ׄc�{�9_�1�r1Xo(��y����87�` ɨu�q��;�-�K��u��U�,s�Dx�x��^r��H��ٖ��fE�Y/8r��w6`�Vnd[����[(���e�	��^��}ɫl��F2��x�k|���=��y0o���9�nd��v�Fa��r�;c�Ы3@��ѽ�5�k,&��&�e���,-6�ɋ(l���_$�K	���Yo���e�=���F6>`%�g���/�>�a�e(�b���Mg�06[y�p��������� 
+��2���������v��N��/� �n�,q"���ΰIL��Ha��59�P�{le��$��leٴ�(u`�I3f�K�*<� ��t�2���iN����I�[i.<�:�aj�-�#=l�P��?]� ^ 渭p���Jp]��S��o�z�C�=�nM���B�[+D��LJ�?xHk�C=�
)'~`h6&��6�bF�4v�Od_x"�M=7`���A1f�@Ő"d��=���<m�PZގj��G�-��֤��\ٚ��JdZ2��c7�:�LS�#��?������o��{��T�lE�s����uB�����̵�A�!ߛ)#Z!���)�[;A�>�N����ͭ!,�t� �J��#��F�>ǎFm�	�����t�ճ��e�x-��NVް���~	����O�Kk$T��͎�F4�Ԃ'qP��w)�ƌ~`܄�z��,z�iS���߀�.�oHCw�:���q�)���:�{��K���E�})�@�U�b�f��m�tP�����)�X�F8�nAӽ5�0/�x��78B�~.�B��tUi��|d9Ł����k�T�zt��O<��F�qz�j�4�L����<T܊�A���@w��Sb�򴄜e�L��96f�Z[�����h�?j�yG�}x0/���?K/�>�����S��˴�A��*�{-	��>(����N!R����;�b�k�	@�EX�q�z>��E[���%�UŚ������+��5��,aa�/�H��+8-�U{7�@���^�6�%���4�>=i���GJ���=?ɲ��#uEY�B|s��3B��d�(!���^;��l0���s!o�z�; ��0����T4i������B0�Rv<�K�`��8��@�	��|;&���2��bM��J��p�ٗ���a��I�p>�盓6�ܞr���ZIW�e���-�3����׌ *z��2ͭ�$���5 X;���`Y��
���Q�6�$������:f+��\����b� @�eM�I�:��!%���3�~�R�|�	nv���e	�mc:ժ�,ݿ޹��l�>�7��~��M5�����B����l�m{���-�,��
���e+�
�aH���U�@+Nݱ � t�;5	A�E�M��qG)@O�3@������J)�dS�bo`�ݷ{"���}ȻDA�P���.��z����l�H�u���,�<����RD���m+�����,�Z��B�֖��Rh"ɼW\��(��%���7?�S�绳��!/i��٠�i�S�s����&5%-��W�7�����Vק_��R�Ϝ^:��l
�e�ށ���Ig~4d�q�n�j���J+���(�D�}�w���z ����Dnl�\tD���qV=oک�f̂1������Kr�q�uH؆��9�6�bC��<K�qb���Y�?�B�x
�Z�U�5k���1� ��{`�b�i�'�0�ק��� �-�=��A��~�+�hM�9�9��><�0�\��{�E��Ż�C���;q�;Au)1���i���5�p�GV'�-r��ª��Bݍ	r�/�,�_���[r��� �@��;/"rTG��*����!�)a@��G�Xƪ���)s)5
/U;h�Q�P@C���g����l��3&��S����f�;Fǟ��y��O�"�xJ���fghw������7�.�$�hNv̄C̜��Mq�w��x��Ѥ�}]���z�ٙ|����:�LSNuF�8�H�B<��#D���lQ��uT��HyQPГ�Np�ʂ��` ^@���#���y��T1��6��������m´�1ˀ!����~8>Wmg�5�$R�a�X���e��ٴ/Ke"���7�w����\"$��R��I�ƭ
�>a-m��L�ӫ4>hA+��w�5���U^��D�{�핕;�tr�v^�_&L������L��摎�f��M�{�D9"�1�dM����L���r$�3��1�Ef�B�/��F&�T�"胩	�����P�d���\gH�A�;\Uٕ�O~S��M�0��(�9�RVF�N������(L����ڈ@r}�N�[PK�|�RC�;�s��,�1j�c�����S�ݧ�&�W�ѷ�Z �-����)�.G��-�Y�����xk_�Z�݅����?5w/��&9']B��J�hZܻ���<���̑X-
�?�+;$��.r_�^�)
F½���n�i<��%���j�'�X.;��x(UH�������0�'2$��q��'��-�'m�j�ۭm��Pf�� �3���"��iNMRu�1)�\R"�������5�6���C8dF�� ��'	{��"��'Dpy?�ˣrF�U�����t��<@8�vD_���5~;�37R`I��L���"�֖���_����x9ш#N�T�R��i�}�8�>��,c����:���w�{T��_��%rb����+򮮣���'V��S���GFn
6��,��$m��ž4�O�@��i������RcڰUȋ��������G�B���R�;ó��D���t*��r�L�޶���� T���N�Swӣ��&�T�y�	�T�&�e�v^Y�j��W�������f�];O��>�d��_�O�ߓ���G���D��7�\)q����@s�rG�{ox��+(ˁ����p�c���+G���b�9<�-�� >t���7���f?�����f4�!��e���\�uq����4�W,tb$��r���Sy*A�2"��pq��T���q����%O�k���i�.+��%����'�{ֹ��v�H�I#�{s�\�\<�J�(�J��"`�pI�D�.D�|U�y����:4�����p�ɉ1�n~�8��r�f���c �������� J-�'���c��Um[	:�/�XG,Z��K��g)M�j?�vb7����C:c�	�
ߊ����%`g���Xɚ ��.���!�	!qq{�o�XqGԋ�����Q�\��W�;���<x��#�x S�q���B��"Cx:#������a0>3�FfcYO�`�:R�;����자�<�aA2&�m8�
<(V�j�����-�b�Jc	[+o=�C<Ĕ#Fy����Bc�ܓ����4i�-�yK!Ѝ+]�^R��|��#8�c��pTw��Lw�y���l#��P���W�n�"$~��0«�|�#���� ��1@�k#+��9�
�UR$3r���$��aq ZO0o�A#�
f�mݑ��E��Ы��l 0��=�N�H8��;�A�sVĿx��!E��r��3!e�#czf���<��I���@�_��?pe�D� �&>�!�G��	�_��%L�y9�!A"��mQ��^z/��+Ø�|U��JU��y	Ŏ�����I}K@Ez}Ɍ�����2�fL1@s�(�=_\�, �	�er��/�$�ڝ8[8;1�]���߮Ǌv�I#��	l�}�d����&|�
�^�k��)ɗ��t���hb�K%(g�Л�<y���mO�()�m��t�c �/�vj��ɮ�R���7n���h���	��A<���N��di�c�Ϳɞ��Yg��ZOGO���~��� �wo �B��%V��k^���$�j�aϴ|���0F�	��9��z�t�e ��Q��w�z�J��W�?��G.q^-�Jq\��'�&��~c��&�<�{�g�]�Z�%�u�Ƞ��o�3=%�ce+�5���/5�� }�D�.~���ob�����n����/(�#�V,6�L��h|��RAsԅ�x���A��l�4��1�[;���a.̤���^'N6��1+U(�S���V�\��o�ֽ�i1���$xA
.��T9�Y��V+��	7	f=�� �n
�W������k�j?rAzH@!�e�x����IGܑk� ��^.@t�ª��>j�O��wm�P^X���L��'5�K8�l	�:/0b�����뒻a��1.���	���D9�LХ䤚�6��N'%UZG���~�^
�1��1�*/U�wZ{p$�ܤ� E�')�K�D�,���X<�[$����|ׅ�^4K�����������w����5���	���[�0VN�ǵw��ro�����.z��?	-�V	}n���@���M~���kƛ7c,�;ixd����W1; <�tp����n!C<>I�)��5h�����2O��>#@��S'sc�*��F�2�����,�l[VYY��V�}���my��E~ۄs�̸��Һ6����U�b-9a#�Z�G�xH�����@4$�Yނ��]_Κ�[��e�cQ��g�����Y�[l�i���sȹ�*_�f��P����α�oM�1���]?,���mK�p��=�	f�g�!�x]P
�1�0I���Z�e��Vǒ��>�;A4�}?�VF�].^5%�O���������`s���6HU
�����B1���s2����e�ޘ����bm�������dԽ��']��� ����,zpSO��zqB'DY[5�G� �8[�])�xw�z�P]A��H��ػ@�NN���H%S#�r+�f��}�}P�����������1�}�X&�0���w��Cq��Kw�q�u�&UH��+���`j���A���,/3�ih�#�Ɉ���fS��َ��)�u��"����_���*�������黥���o�8��z���Q �,d���p�}�
�nwڒ��h�c)�b���5�<��E0Ku�S ]��+����S"> &|��H�W��qVe9O�a�Zor3�c���4	a=X:v�1�6#��x3({5�_9�AdX,��6n6�����B�ې������r��mR������fJl��VOu�6��k �?��z]0�G<��4U���9��a�R��_��ԭSni�[�$���TReg^�@J�b�L�����W�����,�;����F��� ���̖�L���a��E�#1ki1<S��w����,3�8 B_��Go]�I�����j�8m�&]E��ŗV�/���������kш	pAe����E{v�R Y�����!��G)�hۖ�2��!���@�PG1ac�0yEZ�E;��UH^0#�W��+Q6!!�������_��M�5��7 6�@��k
�2Ѽ�:�a��_��0k��/g��|���ؘ���U�6rU)[��ig� Q7XE���V��h�@J프��6��/�_�%4w�H>�6��vh��p�w_ua.�y��n����ۺ�>�̊����ҹ��
�)�"64P�� i"��譇K����E�8Q"�˳��<�I�)�uܫ	�ǥiA���OҚR��qW�r��'dQ��1'Đ:�պ�r��v�:��WLL�'���ӭ�~`���/-��k����X/��:	J0�4Um�\r�{�!�Cϼi�:��ވA�:T�U ��_o��+�;�����U9��bdȸ�V�ɘ�%�S��.�f�- �={��CH�ܿ_ 4v�D� ̛]C����ߍiXg��KW]��I��*��!Bi�4j�Ł�%H%�s�׹ ���,8�5զj;�T���/�,���F(�u�C��`aa9@��(��*�rW���+2��>;A���<Øhh8�!�������(4})�<��T��o�o�}�c��?��o�vD$9������z4���i9�.8r�������\A���`Ȫ��+o���q���2!������|U�Ӟ�*i��)�~� �]��T�0S�6�7�^�d����3��e�1/DW3��X�,���/.����"R��m]3�)A�O��O�T��CV�W�o��aV���7W�N-�x��HN�z��=���%=ZA�H��7��/���jD\j�K�>+v�G��`���Q��+��%}ڛ_��zJ�=�B>�[���ɗN���1�9.����ޠ��@5� �>�~F|HZ7J��˾��mQA�(��J���?��.	^�i��n�#ۘ_��1�������˜��Ds�\�1
�h�'~��.���[�۔�֟��er7�C�����M�i_���(���[~��!G�7mf��A�G�QE\����˲n��ԏY@�����s�L�h�qH���\yR�	��!%��!��j�>���Sn��]��z���cX����llI�xk�\���$w�ZLv&���Ί+8�P�$$sy4�����i��MB@����Ak��{��q&��6����,�O��=��LC��<�rP�_��˾~��K��]��G�I_�S�u��f����KRw��G�Ϲ�����o<���8O�wT��J�+<L����`���p%��l蟐� '[j���I?�"3_����N�fd��Qrɝߕ L�a)�x<̤��4]��}�Vm�^H�}9��PP�;�@�=W��ͬ�t���N��ho]��dAEz*�j�_�=���1�u�»�v���\���a{h~5Jn��M`N��)I�'*��I���_�K��m�$�5|��L͍n?4���'�屮l���o̷)�Q���U�Dx�f�o��,�'5y)������Zz=8-�*�1|Ѝ����Ҁ�����wG���f��K��7O6ڛo?�<ź"];�֐'�::s��������"`:��%{�QA��k��M����O'�`{�CfL�1n����&�F;}
����*6">��+��󵵗m*7vN��;����W�p�B����a�L�����qz�]����gv�Wkps�7=C���}��@�'�h�Ì8�3GH]H�[�;��V_�	1Hة�"�� :Y��7xB�k�?�������9J�a`^4�F];�2��4m��-[�覃lG<�}$VF3�u��8�p�T��wg���~V6�h�Fљ��H���D�|����`yG������2Z�GP,rNVnU^mDv߼GS�R�d�d)Z�Y�n�%Q.o�^=�p�V$��KȄ�1�@k�TU\IK��zᛳ�p����M����0͸�;��aG�����gp����[���Z��	/��X���6�9	���->�r�=aYvJ�G�?���71�K�©xgx����R Eykm�����9.���l��~S�}��.�6FC�w�ۚ�©z�>����I��(��|�x�¦(��~q�����gRإ}��g2�x��F/ ��Ԁ�z>�Ǵ�:Q��/�q7�S�Pf�$\��ݘ
C��>�+������,�f��K�櫳c��4T�/#�.����7m�%]��wo9����t�d��{Ld����"a[��Z��/J<F\N�麈-J�&3Fq޻����=Ls�\f6{�b�k ��n����gم���]/��b��~I�"?��H�s3���@@C��q�D��X!��o/Ց���pڬ��u^�#Ȁ��xCk�r���0_ܰ�=�5f`ziMH�t����%���
l��i�1Y�`� 09(�tm�oB�Gq4�
� [vk��Ұ�d��Ꚍ��ᤐ
���'G~1[�Ř@���;,/���*��ߨ���/��b��8i\���us)����y�8���HG�D�<�bje��E � �|��f�b�Q{�ߍ\�
�ʇ�K�d������H�~�u�)Ӛ~Q��b�!��_�x����Y�݉8W�Gqߵc���:��Ӣ>���E�;�|�>�J���IA���a�� ���PV�w��
���@�A��#��l��V�0���B��A�T�%��o��A
�����Ϩ��ٮV�Z�r�Q���Z�O	k%��ȓ�qa����bV:Ġʶ��	���:��D�q��g���-��/��쿥��)�N��J��o���)1a{@�[Щ�p�6���
�Y��x�d
o�E����� ��@w�,����P�ʍq�Uc��4b6�}��7v/���l���O�(g�ً���g�ݜ��M���)3�?��D'�0U��Wl�CdiRf_é �1�c����F���h�[���:�&؎>�#$���8�i�b�bN67juX?�H{�r�o�[��u�悖{������w
��V��(�ߕ2�c�R>�ȹ-�7�a����+)���������J��"�$��q%�p��4=�L�0�;�2�>	VOL�U�x,)��fJ�0�s�DA��r�hQ��6����8�RZue"10Ǡ����� Xyi�7�?݌1R��^v���Ϥ���I����������Nޮ�"���j+aE(�k��߸U�u��i��H.���%-���ZÉ�7���x�J?�`57���vFv��4=|��¿�f�d��6��AS���"f��'�b�G��>���U��@j�wP����'HH*��f�Տ�Nf'N�FNy
p0�oȽu�¡���Cy�?:��YI>z,�Y�iLZ��A�ل_�aX���1Z�έp^/�Ip�/������έj
�I(�����0(oi�:|Z7g����%�?��Ѕ�Y��9��	�	.YJ��Ƃf@�I9�If��P$'��~o��n�N����ܛ=��ll�˳�/c��D��֚a���4�C%F���/b�~wE�5������:L�GoiN�$��"������ld ��@��dXa�0\�V����sɌ�6�,$G�D�g�w��|f�u��Ǭ�mr�K],3����c�$�Ӗ�c�1P��(y�V��[x�䁱m ���\<}�(0E���*ǴK��,IB�-�|`�t�O$ ����$�2E����}Њ��a��1<m�>?��7��-��"6�P\�d�����3�I�?�)�$�@��� rq�)�H��J�ǐ�Q�)��7mJ�����3�����!o��rZI���-;"�N��,*��x��^�޶<|B�a����5��G�y�9�g�'O?Z;D2�$I�^7��Ƀ�3�SX��Ͱ]�w����6Q�o��s�zW�����g,8N� ��":�-�2<j\!.���� D��DN��_���^n�NcZڧѦ�[��CC��j��!Kjl/��"塇����,{��(�P��"w��B��p�e�q�k!3���KUz���AlP��ܛ�R�8I��x��m}�d�'�>~��CD?xt�L�s�\����/"P�I�*�K��0v�$��>�N�S/<l����ԍܫ=[�$�A��M�ߴ��
+�V%��xa��üY�&˶j����:�b@�UX��r��Sl�V�N)��{�3��;L�;�U����D讧
RQ?)Lj�/����W�4v���i��^�qt��+5��e�)����4�P��N�u�!.`���B��u��ς��j}�� ��1�b�D��
_v�ۯ��]��<׬4X�����ƀuH7�h P���h\.{����/m�O��v������'��~�ez����!XЬ�OH�J4��&D��p��Q���o�J��E*�V����������g��m������<q�zAi8�&������
�8�a.����� !�����0x�tFlL��p�A�r(��o�-�&�N���=�"A�(�~a�c1���mBێ��Qb���= �Y�������Ck^^2;LI�͉k������(��ؙ䤨���-���9�d�<㱿�m��9^@��ݨ�!�!Ԅi�1�ˠ����<�k�ه���Q��ﻭ�,�k���3,��ħ;O+t��4S�H��!]��gU���D~����X�~P������۲SV�Zo���v6��_%�O��Ka!j����!HP����ud���3�r�\���p�2w�+;�4�;b���X���n��!��#]��m�� ء)�(ڛ��ȸ�z#�D_q����*CP:�V%o�9E�otBD?߯�[_tC��ا�@w��h��FW�p9:[��>���whl|��H�6���ˑ�l�w��`�=:2���V��Н���c�Ob
ݓi[�g2��[X��g���8 fl�sg�;K<�p�,�~k|�.	Qg*%�|�%���-F�LDۃW���ǈS���EK��9P��3L"RAWzo^|j7��/%��M��ޟ��RX�?[�0 ם�a���(�I��+�5��8���ҡc:�@G�yy��� Gzr�w��y�{S~���ﶄs�F9�\��㝽Q7�%��d[�B(l�=�� �Ec�\��S0ϥ$����F.�rm��CO���x�A��QG�f�kT9.48*O��};�}wphN:����%&)������^;��xHj;JMX�	������b2q��{S��+����_9_&�x��U�����)���o������y��*G�� a��%��(k�ȣ�s��Y'�YP��1���Њӌ���''��R�m/�JO`*zt"<�Cj'�y��u�xk������H�R�#p=f����1�K8U�V�qˡ�1*(
�#�����(�tYBX��'K/A�Չ��3�i,C�#�;sx�l��[��]���@sK�,��/�.j=���v�e]M�<C7Ik�|��ɲ�,[�"X4����V󁍏A���w�^$KV�ر/=ZҢ%-P`�P�Z�I<w�Nzv�~�@v?�Ҿ�s���ζ�LN_����,6�#�����I�8n���L-�O��#<w|!:2�F@��;De4�3�����.d�2`�?k���<���bX�$���{N$7DIM�x���W����/A�PB�A�1��R�#�r8�� q�7-Gkt�(����n��+�#dɆ�q�ʒ%3|�M�E����ƕ��!!��:��ra
�z��G���v3� ��w$��lU>�? 'y�V�ac>,=�6�ۼZ9	(���p+���<F0�I��%��@M���+���CbvQ3�7������j
���_4�Ku�x��5?�}6K���LuG�jDu����s-C�ݤ�~�� �ʄC�gE$PnΰS˂�����c3��Ӌ���RW̑M�e���u���bC�m��a{.���_��BmL`Q��v$z7���O��%��/�k#z�����%%Lk����6rĀTd+6�~�ܐ�x.�.�e�� ���%t~���,˘j�*Cl�/���t�����B����ܦ�;�� D������ 8 ����ayhH�@M��y i뺲�������Dc��E�o�yРRcL��S_f.t�T��&2����>U������C*J?3��~;ԐZ�U�\Լ�f�_��lo^sd�,4�~d���FN&���.ɅE�#=�;(t~n{�g��#if��95���T�&�W�&�
sP���F��\�- ::n�$�}#j��`s-��l]���Z��?��B)��Q��bMЕ�3��O'��"xh�v��ӠB�b�F)%��������΂V4�ٸi�p����+]�-}b�D"�w3%%d����v�E��������&��,\���r�=-hk�E:;,L�E�P3VQ���#3���ˋ�vٴM����D}�#_`����X�����)��IO&�hWXr��@5Bi�������a gy*�b��DY����m�v:�a�� ܸ����9Y%��N!G1G;�5���y�U�T��D�����p���;<��w�m_#�	A��8�	ݪ�芅ou<��|}��K��
�͢k�Z�
T#�-
��{�B�F;.p����������J�r):6�*�[����q2.���Z���l�j��s����x��;-����Z��,����`��
�<����5������D
^�"	����u�����0Ļ�K��.�6˗�@e7���1|�,�'`�z7Џ���s�DV���A����%��ʨ�8���o4�3H�^_L��" n*�a�TkAM{��y^���5u�f҃�r����%R��ci�aC��hŪ�!�}�����=���Fޣ,�G	���U��w���B��������ز`�{�,���?�D������b��:��Aꍪ�(��\({0����'���r���/�[�{�A���_Bc��g�g���īp^�4T�k�.�?!k�Ik{�����G�U:�ܿ{�I��="�5������q�hė}�?Dn}�y|��`�������F�/�9:P�c�(���}��`7���;������2�������d�`
Q<�ɱbt�z������},�����,����"a���l7\kCi���d ݥ�UE�����p\��1�"��J �Yǫ�(M���Tz/�A���
D�Z{�Dl�y	 v^T5  ��������_��\[�ܚW���q�*��;��ʧ�'�=�ݽ�qʃQ�Ƈ�) *f'��Ǡ�3��x�#.+,i��?V:�U�u)��p=���>�
��g&.�ׄ���h)@�:z��M��M�fn�-�� �n��q�T
g�6�X \�ߏW̼�X?�����b�5�2R�Z��sKv7�7჆	]8�j���C)%����4qn���Zr#�4lp�wd���<��v��I�ͶL1�/�� �Xd2��NH .PI@����mWI��R$�2�)rIF��8y�I豘=l>��Z窓����ڍ���(qZ�ib.i�ܯǿ�U�!��Q^� �˛�H'Z����H�1j��6�^س9��Oҷ!�Զ�����z�gr��q��T';|�E���\�T$)����	�O:���U��8�Y���9x�mCA[���yJ[=��**�}����$b>�=�Z3�o;,��!SeZ.k$w���$!�pY����>�s�J�~�������%BX�?9��Cn��*6��F�%n��v�o@�c �>;��[�!@[�o�h���k��%��>VL"I���$��!��Ы�Jdo)�Y7�8uG��K3�����D��H��|�|�|0�
r5����?I����M��meG6���l�ީ=
A��L��� (0B_͹�S�˩���-�Y�3�4��`��T�fh[\%(ҷajT�yvfb�햖Y��Z�OE|yF���9�)C!<RjĎ( MI�.��k^�W}b�����y����+����_���?�Ah��L
S�m�z�q�J��z��D����\YQ$@�؊�w3f��N��A�D�$�n](���Ѹ�8^ {��-GNPNViΰ�F��M;�ymL q�p����ܿ�l6�����+���Hh
!hJ朅ݎOH�\�7��מk�5�9hs)��$n��tA�����x)(U�]Js��q�b�A�d�������?�H�,��i���� K��T������lJ�z/7	в�TU�w�Ŭ?h����O)�x��VYS6�����o���/��%�����G@��'�G�Ճ�S���'�g�QT�\����J/�i��L`��_��l���5�]�AX`��iH"�(f7ś �э��2@`̲zz�b� /~�Cs�:�n���x�ZF�Rs�Oa�tZGF����@�����(���j�n^�k9qT�ܜYs�+DK��m@��Vt8+�c3�l�0��Qվ��1������.��6f:b	����Ђ�D�e7XX�ː.��x �B��Ͷ*%��,onX�c�IkX����f�*x1��0>�
�IG�>���'�x�1!S8X/k��L����2�כ)B�m�~.���;?��*i��q�6X�K�*��N1�%Oϩ�?���������q�PA���%���(ֿ�x܉�<��Ař�1�O�=�fݠ#e�
=|����-w��s}����-��lJ<H�X��[��,z��4��)��S���2t(�����v��`�ɘ`&��-
���6>��KY��#v�ǣHB�aPY��7��12M�	�Aw�c����.}b�c�2#����<d�����{��~ZY�;aa(�Ftg	.k@i*�~j�U�#�XX��1wMR|i�mH��}��cJ��T2]�i`XV�R�'c��E��V]�}b�fl#�4���~����a���}L����ӈ� ���O��T���]� ������#��Di� <�#w-�_7S?�y�I��%��_��>���=:���b�PL�Y:iPnWf�l_U�x�(ij�wI�F����Ӄf6Nq|����x9�����rǈ�"��0$:$[}	`<��������Cߎ;�5S�U���-!�܎�p��^aĆ� {{��Ԙ`�N��A};�=�Y��<w��|��4��(+L�Dh���s_�֝���D(oV������;�C�XQ�a�[{&��De\��޶q@Ve)� �� ��m�*Ea�f�ɺf��i#�[$�f�K�l�vi���sUSe���XIx�{}b,Ak��3����xR����+x���?.,�zv�d�͠t؁r���c�,��WӸlb�d2x�Q��[_ 3y.\����Y�3܏��	� �GIHX��2z��4�/-�?�Al����b$�2@�gJ����o*��^K��ґ�{�'�Uz=�`��x�(�;@��
J�ʣ����(+��X<��täQ�� ��YԚf-�����6�m�Nfbw����ۘ*�X�x"����݅�ޖ�%08�qVRBF.�� /l\r��m���~��Z4�#F;롡꾖)�s�C4w�Oԕ�����۹�3t_%D�(Dk�]7ч��U�p��"�qpz���5q5`�{�&9�Y�u`�MP#u��Y�x��<�M#,7_a���tVt%4Ŝ�O���qB��Ũ�d�ei/�L%4�,�*���嵽dDƐ��)����sTC,�a�O�J�L�o���F#�����.�C�]�<�˟h�{��^ݩ��3��%(��V��9���`�+�C���7��Z�Z(��?
��A��ء�\��r��B��F�_�Ϫ1=�I�v��� [*�d�LJ$ml��v:3�a*��8:��(�'���SV@;4�	��	 ֓R{[��7���SY�e�����'ۧ6F��+w�_��+� ?B���k��$l�*N�1b��� oMc���(X�� T��`n�U��ǿJ?[WvGEeu�F�װ�>����xbg5	\uu ��i��~Qt"��-������4CL�q���\���;��U����h��Y�>Vn�ߜ��]��R@أW��\��$q����&� �G��+�WNyI��ю�5[jrۖ:���#����[�G�G'�|�g�Wy�;�RP��q}���mZ�>�Au�ɛ�6'�l�}J����xAN�訏���56��O�tI��6�v�wI���?�fV�wDք���{NQ�GUZ:p�k�t�nu����j8���T�Y��.-$9��f(�v��(͔�5�vh�R]ΐw����2�!03Ù;a��z��i!?�<d]d�y]���},WD ��჎�U0/��i�4O�~-�a��~�KM�p�t.�ux�r���`�M�j��|,�\b�Ef���K���#4���i����Hz?#�8�c�:v�@D�*��M�nmq&�m�~�	A;'>��	�I�w����w������Nf�w����۴? f�|+�����NW��k��1���$Zo��X��5s:�|m":�LDԎ���v>v��i�Wz��
uv�s�'��"gu�<c�~Br��DJ_@�j^�Cc�?ֽ�C`^V��D�Ip�#�C]E�+^��c���m�R������N��A�,����DM��Yz�A��dPG	_>��Rr�?�\����c�2�%�����̽�NJx/��h�NT�8��徳��N �[<���(;y���Z����̨@���[���N|��$�cos�%e�U�g�JwEݫI�\f�i�h/৤��	��`�"k�G.�VF-2ߝ��h��n�/�A��K�k��{2Xt@����Szm�����u*�3t}��_�~�tV�%xO��d��䇭��X��1������K$�4�\}���B2N�1�/�Pd����yH��Ы�ݐ�k�`�5^R���av��ez56��c��&i��5)�n7�L�~=����tj6Y8|#4*^��4����"��*'����:�#nK����3{ϸ�&�
<�_rq��7�[�Ü��	�}9��b5̹,q�v3�䅈F�H�W�k���a;�c�06�u[ku���ᛟ@z�!��t���j`#�X��f��2 r(A������ˣ��1�,��P��n��֞�7��|�O�7(���ļ��*��n\�&<Zwi�i�S�R�J��A~ѝ9�M7rE'��o��h����!�+�6ſDjW���WD��5�OX��٩-�Fr$����I{v����7*��E��1,CY�V5�O����I���a����X��ؐ�aM\S�B�L.��k8b�%Am�ZS�<w�5���-JgK����q�x*H���D. |�ׁ8�l��l�;^!1l�J�eFG�Yo�'��Wof�E�t���V`=m�dP�!*���2aq�`ǶzT�C�f����䮿�E[�m�c3�_��.)@=���_�2��;Y^�`jg�`�B��.�?G���@!�����1U�{\�U�������}��(��4���l����o�F+��7��Ai
'xb
�5|��#���7�v���<�+��I�D�װx���ԅ�¾��(���P|��}j�DVĿ��{! H+c�<C�C5���C�̑�Mab+7�^laSe���>�!�c�ngo�������� �*�)sd��o�;�j�A8�9[��(_Y5Z�4>���%��3�6�Te������S�/K�K�V�+��P�������)�,�@:������Ⱥ��[
���&�U�UO]�W(>1�z"��\K*�SS�Ji��;T��� ��1y�r�����)P�
˓?72�rZ��W B �U'4d�0���|7 �%~���<���v�Uo���d��\!��	R!�h�j6L»�'w����CvV:���Ĺ3e#	�O��໖%�9fU�B��o�`���oT����R�5�ֽ ��I>ى&�~2T�܍�	2u-r>�D�g{7����W���
�_�;��y4n	��\��v#�J��;U���\�t��ȝ����AO�ێvx�ZP�)rw��<��E�x^�+ڍY�j�ன��T%���z�+_E��u�������wغ���[6t?���G�<�c�edK�:}�=W��b�h�(��%�ӝ˹�IьJ��f1Oؓ�C ��#~�p�bB��:��%I�1ܪŀ���ƭ@\'/ekBQni���Z�E�?G_9h�i��α��|�i3?JDk�B��T׵EW��শ�MͲ+w����H,��W���5Y�>�L#��,nw�2�_ƥ�"�nٷlM�^�Q���:�:{��)njw���y��<���.��d9�|:4u�lp��տU�O�����U�xf�9E͐��v�T�oH&\L&�eE�).�{�!_�$ݖg,oFP��'�qX�x}uռZ���'��l�P?�y�>x��܈����Slj����4 ��բ�MD؏�A�m�-��g	_��y��������S֭'��������z@ 1%�r�sN_Ϝly|�$*(B��E��Z�����O������O�6�V(��-)ؚ���"������է�Rk�kc����2�^^s�mZ�N�)���k���3e��?/a_��S\UFc�}����(�����/d�ηa��֛�ؠ�qR���"6n��)���]�丨��*����e�"e�m�5>��k��
ٻ���ހ;m5[2b��t�Lږe'�F�]�|nR����e13�,��Z�%�/��~���k7E���e=V�����y]UJW�B �{*5Gʆ�&��j���}�Fw�jS@�W�q�d����q�G���E�Y�\!P�pgnC�� �h��_b@^*!Ӯ�A�cT�6�	l�G�^M8Y_��NC���^��@l��:�#��k�$���;��^�jF	�����ފ��ANe�D?!Y~�9���-�(��5|�A$!Ү$r/cr�%��)�;�g]��h�f}��,�mT_�BlC <�+�'.�|F��d��Rn�Ⱦs�`C@� WB�����K�\��X�0��Nf�m^���ܞI�1���$�z������`�b�uq!�|t��,dx������6P-�_��&M�ǪN��-�}<�@�ύ(����cc=חnp�0˖�C/�d���4R]�7[d�|G���sx�;���j�{6&5��:�	��m��A�,5����?E�D;?�̮�����҈=��
D����&�*;X�6Fź�P��$⭁*ώr��҃l��j��}����$�)���iD�W��:ط�Ԁ�A/R]o'�˼UO�76�����\�M!c<n�j� �r��L?�6�?U2u&�`D{��ߵĢpZi�B�8��2�9�o�7�X��j2��WEA˳YBe������-Y�T��J,"r��`!N��Nk^�^��L��w�*V}�!���VL���{y��qv�N%�J����L�����ވ��pvlQ[6#H�~F`,�d���&�X���>[����f�ǽ���UxD��V�S���!�-�5ᔌ< ��[aƎ��;%?����I��b8|l�k�$�|}7���Jb��^�̓0Y�v��2�����ZqeM�O���	�!M��,�B��a����� ���f�I��'\?7���tK��T�I���^��E���8�7�b�)�2U��*� ���u���Sf�-�o�s��<�lJ6z�Ů �x��>T_fi�N.��j���V��C �m��a�7j���Լ�F���XH�Y�'�hЃ���E�N�\~��:��j=J�<P��V�P6-|����"�b��4�m#?��2�Җ�%�:�
��,����)��rv.�
+��NqlI�r������vZl���
i��S.�W���Ƽ����@�Wdp��oy b�5-�9��tc]^����6CK���c�P��������?�W�(�tG��i1��^H��c� �	Y���Xn���r���#5H�כ��C �;)^b:O���M��w�fՠ=Xn7T���e���8�6&n\��m�7r�}h@��jLG��G-~�h1OJ
P;�{-�nax�t��'l����J��t��{�u]�z��|c����&J�>)�	�|$%�<���ݤ��:��Lx(aBڱT��ĵ���a��M�qӋ5u^���Km�s��SS������۝�0#��J���ꨁSvh���R��<v�C�;���Ԥ1�Yꉅ����ޥ��)��x 9�XNHzZɈ�j>�c%h`Μ�x$�≀&�����|xP�F��ϼp��Y�޾�DڄO�e��۵�i��������������v��\�<yY���|O���xy}5�����x!λ���	t��f,�uvn�07���+�����f�zX�CVkN4� \4P&�EH�^y<*�Pj�J�����%!��*~�tbe���0���,��~��Rm�\�'@B�`�5T�M��a��Q��kS T���H�6���M-���Q�r���a����Y(����f��ʪCֽʐ�g�٬��A�# @���1�s�a,�p�%�����ta�y�NC�\�b�l����ؕw��' ]��
-Bq�o؏9��K�Zu&��*�a�}�ga^���2��n�)[gl�������nH��S��S�6���Vs]u��)6��tAR��yfM}3���ǥ�B�� �o�� �`���8����}�����\�N'vv,��xK6�Z���b�vf���D�0��E�����$�o@�:��s��E��F�P�LA"ƀ\%X)�QkPx�#�
/����w��m���'���,�)Ǻ�'�����w�mU���#^��QT������r�(�_�J���B���D+�\��?�%������R�="bUSSi0wj2zÞUl�W�T{M}ڱ�㠵�q��e�PN���t��#�7�Sk�p����Y3��!jQ��?l
+oˬ0A�.+�*p���.��p"|\?�=���Q����~�2J9t��ZG�\��jEZ'J���ȑ7�����(q���2�U�]9��z��nA�k
�w�6�'����'�6��/RO�.}�0�4�9-�Y��h{�me ���q8ۖ�q�AK��W�K{�8�s��ߣ�,�w"�K���0ˇ�j�.Q;�3�~��Z�p7;��oLmw�$�5�s�w�
���9��E��ѝ	R��	kg?ԗ�PO��;�� ���A�;����* �$q��Xb�u�k7���W��a��@��D�/>�E�XPg�x���pȣ� {�L�RST��"��������O��fǗf��K�=S|���!p����
�J�(Ye/�76�6��*õ��f ��21Ym/����X�"؏������:��v]��j�o\i\���Ef��!�z>��L/IPD��oض��CyA����[�^���H��%�ǉ(ҬYE�WɠX�a��XX�OK�H��==�&�[o�硈�}p�kfq��U�%|s;�l.��yFr�M
��`�кh�qլ5���j��.�����s�"�iz2�a�E���B%@k��3�Vh*��YoN�IsRY����)���n���4)I.�Z	;�-@���E}�� 9���j���g����4n���D 0l��}�V/���1�1���W�5Fo)�v��K�.�/F�=��T
�Cs�H��bX*�?X_Ns�0x�4I�7M��H*�q��a��U�����=9�C��me"<�Bq�+>��-��e��T�%,���1�����sEI�,, ��WЖ�
�ع�m~^��뫁�S"�y�����%]�;#o	�`G�ۚp�zC��T���>z��nM熡�9�Ņ��w��@!?�|	�~��ʘ�?���`L���71�:�dRܾ�
X[�9|7�W2,k��ab �t	KgZ���g�X�4"ˡ�z
~w��(z��� 5�4��	��R$pގa+*��wk��������Ԥv�k�R%\����U:��2hL��Ç��i�us/vl"��5�2���9~%V�r�l~!������~��o�����	�1��WO�Zk��V����U��$%B.QPcBM{���h�UO��3+veʳ��>�q&Vt�)*��B4p����v�D�uƫt�ڑ�Vk��<��]^�>#H�-�*e��;jW�7l����4�92�筀v@��"3K;O/Ɩ��ve�^�0�k����*�:ZoiB�h�J"Z��~���������>�WB�y)ċ@�Pݍ ��@���4Ҝ0�r�G�d�/��G:eB��nC���˄�l��$���#��yx�f��U��s�ԧOp6�޼i9:8Z8 Zғw3�������-�aϻu�9Z�H�;�2���qCʚ=Ŏʯ$ LU%d���l��D���{}Yd{B#�BCQ#?���x&��ҍ�Z�U�{[r�s��Ǥ�~�����z^$g�*��0p����Tt��|\��P�j��N�	b��5���������y~��H��r�73��o��.3P�N���ȫm� �~������J9݈J�0w]�2מ,�2G
��V�5 ���n���]���9���T��sO$�����eo�F��N��� �0�U�ś�J����$��W�o�����䗘v!��ꒄ�;�u*W���d~��*H'pc�]���O�Ls��mms������h���g��q�I)T9���^
F�.�#�ꫣ��ڀ��[�aV��1�m��7*�A/��`������K�S��j�M&JW������X����Hqj��%����Ge���*�r���A��Ll��鮤�P ��N�q��Ƭ�
C�l����i����\�֩�� ���R��R���r)�c�E��:E���.]��-���&�!��g��:^G�<-+(c!;��C-�3O;o�"쯘6���,��SH��ξ����D�з��m9xx����@j ��D{OV��v��3(�bώ�V	�(�ض�҉ǡz���P���$��Z�7��P95�+�{Xc�D�3�s���B>Tfl��®^?���I(x����3���h&ӛ5�_Â�Z�-h�%�ެU�1���^T*G��R�Pl"���}�N#74����@(�(3=.�)�,L*Њ���Veh%�0W U�K%����W[r	W�~��Gy��.�y/j��rTeӳ_9� ���	ĞT'�rC�6�� )C���L�'�4Hm�)L}���U�3��e����&����t]N�=M���Y�Pw�-Sc����<\1�H�t:$.���i.����ٟ�N��NU�߷$�hG|t��mB���<[�~��8_����8�)����$��U]����|
"�J�C�TG�`ڧ{��c壏���8����a��#�P,�ц�����Lu']6t�P�=P֪n�2^.:�`3Y /'��$�Xls융���&H����7E��Qs�LX3zd*�!5��2�ehC������V���if���Jo�{��Q�}Z����U��d�ᤜ�kg��7�ab2A�o��Y�jt�ۑF�X$��S�M�f��Α�s^ûrM�T�J����͕�nT%T���ѯ1�;R7�b�}��Μġ�U��(]�r�B����6�!�;j;���N�$�\*��|v���5;�����"�g���r�S�;>����I�c+�Ak}h������u�w�E1�M��ob��;趯�JOیt�;a����xi��լJ)2�M�k>��-�,�sw�bj% ���[�g�[��ᴥ�|UB|!nV|,�'�^�0i�]���Nw��6��`H5�ˬµݮr�*K�X��˦����M�X��g�㡷�
Y�t{J�5�pU�{�@��-��u	{\�q��}Ҩ5=\�s�p؄s���hi��Hɱ�^��c;� �������y���Ɖȷ�����G�����E�v`:�=V���J�py���d����/u��5���a�#�Y;�E%N�Y��d���q!��p7�\��P9�u4��w`�$Q�P'��9V����b~t��{�l>�"�dV}7�*bE��c�+������ɿ�����M�ZJ��9���P�Rp7�l��0u�g��=�n=d����ǳ���іT�W�z]�!���D�O�~w����9�EG�uLȦwj�Gw<}��Z6*�t1��3b��pd
i��x� �����(�޹��� �ZP1�bn�f$�R�樚q��[���R�ޤ4l�#���fcZ P���3cƵs�k���[� � �V��I4Sۈ�1I���L�g(G���'�����ס	מn���|��}�?�����"��0?�{:���r�l�����6�y��<�T����gvs�����E9���vlƮu�ur%_��鋾m!����&�f"�g����Vm4��T	��x���d�J|�>-�*�rΌ6�皴��B#)���#�W�;�����ջ���jա9<���gm,�?�mi��[�Z�3Y��q�D9ۧ�>�W�?�����䦿��א¾4c��<f�>�O�!�Z���+�wa^��Q�8�)W�LӠl�r�(�{����Z`�)u)�\|��76K��p�A��l>�ѥ�����ܰv�cU"��7H�Z��		����&��m�d��x)T]S����x�t���8�VB2\oP�ݕ�|&�>�걕w7E���K����sz+T�p(<o��چr<������Cʶ�yf�l�(���F`��K"M, ��C�M�d�ecwq��]�w�Ȣw���T�eU���������##���9]vB�`�Mc�����W֧O����!ݬ�'��/j���x�Um7t��;%6�f�}��/tR~an�5z.;ŰQ���X�Y��.�sZb]���L�z�����T8�ٙ�b2a���b��DF*v~:����G� 1l�_�D�4��e	�S���7���hv�!�GY����R>տtP��[���d�Ҹ��c�	y
�}"�M?�kdQlsXAz�	f�c���r�dI|� �'Q�z��ڝ?�p�6�!�)�t'q�J9o(��_�C���Q&�t�Ј:����x���[���j?��E#�'cگ������\X[,$�I�6����ʓ���|�]յ �)⛿&��s�|:)�!���Y�ʝ���\�h�P�V�La�`!�t3�~Gx~�a��ʁ��W�+J���������;��M�"�!E	����%�1��7��2塍��#�Ϛ���ɷ5��7�� ��v���[���TDqnlCx��>���qu�ťc���r�D2�$bJD1�8{�<@�N;e�Ut��S���ͥ��z(�~'�%"77p�[�c������)Z�BT΃����s�|�9<����K^S�b���v=��!]��� L�, ��K]CAy��"�P_L]�^�Y�~��\T0�~�]�o��Fvl��aT���g��b(���,E���_%�
�t��u�X���5���d�	�y2O�����Ϲ3��2۾��3K��5P�?2Dn.�o��ݱ(JB�E� ��y�ě&����*ĵG!e��	n���ɞ�4(m��}Y��ls��f�Hz��b��r��ݎ�]W��p�Dd��@���b�KK����T����[xO�$�b�a���P9Eϯ�v�4�=��O��
7�#g� �U�!��x$�C#6%H�5Q-���a.�k�g ���_�:1����D�����V�i�9����/�u�Ҳ�S����A�vש��囩dP	�xK-j�c��6�����&sM��"��eS[���ꅭ&}�i�iX>����uTX�~��\�����gBKD4pn}Ҟ�M�C3�j�$���C��X/*�t
,P^�H��b3���:\���`��F��x!����q���6j֯q�#��A��jD���X�֩��}�@5-]�	���^<��d��P|�J��jS��I%glKP,�ֆ��<���y�P	*q\te&F`\�̟H}�zŬ �C�Vb����0�ș���A�踂YsW�s~���kK�!.���;��e��vFJ��M.�"���� ����{�o�5�^���W�!�o��B��p+�^��
[)͠n�Y/TP4��.2���:PV��U��+D�N/����}�9S|�һ^*�M�n���WR@��q�B�%�����U=\�G��~!�Y��ej�2������6'4�z�0w�"��PeZ�ɐ/5za4 SY�O���
�;r��gk���@�r�^���cL����ah�PK�G�x0�����A�2��m�C.r�`@=)iz��>p����AI��o��7]��}b�������i�73��`>8%�kZ	 �4����2��P��a��u��t�uA?������-�P�v]��ΈL��',b��$VGvi�5�1���.ھW��e��٨Z���������0#Џ��g�a^:�oZ>T2�pY�k��$���i��;Y���a{t�ZB>�@n2��,1�՞:��wg��"D*j�����
$9M��'-M�_�˸�R�Cݽ�l���������1ϋ�M��#r�D^�����Mx��߿��&��pLiM{W2�'���m�'�q`�-V�e>��"��`p�ّ0{�U�|&�>X�����͛��[9Ga��r���);ש��똈�A����"�iT$w.���#(ô�ޑ$g�� v����:�T��#;y!"��S�o��Pd�s��S���G�t9�Wz`�O�	�u�4h�ڌT���.T����h|�(�P��YA֩�
��!�蚐[~މB����r�?�)�`�]�J���7��`$Q��� ��כ���g�fu�M	��27y���Ee��0\O�M�[�+�j��.��/A�{�������أa�B�l9P s��^Z�Wȁ="x��N"�j4��<[����4%af?~T6:c�v�hM6�����Hu���,���F�ȶ�[ؼ�ެmf���$�R��e��s�i$;d��`C�B��3�.*�2)`�U�4̩�zohOA<�n@!U'<�an��T_�6���]�w9T�:�G�p�И���&Y����	��E�Ŧ�6�Q�HSTBMc��'�=�;��{≌J[�ѢN ��?}v�'��ߙ�&u�9a�D/os%�(9�߰��*�K�x����!�M�~M�:��.�0#�i�xu�Н/X�2^iM��D3�#�0
��5{�������,�AV�,p�s&�cۮ��;��!�	ш��M1�E��o��^xd¬���$�O0�^̈���f�����@�O����4A�L����fޗP̺g�M�P�~I�;����5�/����ɨx���V`ol F]9\�õ�?(��;o,����qRj��zi2�Ԣ&4�Qv�?���.
���2�ݜ���g�nш\���oUp�����K��$�����hJS�F�'2��K٫Q�q�>���|0�ƵF,.R�F���J�7�Q�כ��	�.!��D�r�Ф�G�c�M�*��&)u�R�����q���8+�3�j�d(�
:�r��k	#���Q}�cI�)#%��"=oF9��=|�h���ǬD$��#�'�����|�Y��P)_�K�a��K�_^N��l-HZ�����I����1j�:۳�
���pﴉw�[�^��3�}��'ft�����e$��"V�5��WtE�i�~`��b�G���sQ���i3f�@�����7Ą��u���kLeH���2ȹ��&�Nd!w/��ƨ;�qx��/��br�}_F+D���Tx�*���S�["�"�,�҃i�YH��k7-ru�xv��U�QX?:�e��g�I�F�h��t�5c?�<d��ӫ��G#ph���-t��1�HqC�G�A�����O�H�]]��ȿr���t	m\ﭗ[�ҹ�Կq�t 7�s�t��lxu��rzwӭo�G�m����-ާ]�3��ec�	�J�7����/kY�%ޅܣ���xBv���F)�9��<��l-�����K����lC������a�
�!Y	7���o�Tz���sB�a�����)�`a���.��؇؊g:<K�����ǥ����[T9�*�W��KS�.��c���R��a�K��
l������<��{|����d~[���9�+ �(b��U��Bt����3_vm�e-�)C=l
�Qת'F.�tޞ�P��Q��?v�&\��(�rGF*}�����7{����ٍ,�WQ�"P>�����g�nd��y0U�T\�Kr�hD��=��u��������J�-	���7��o��x���]b�3\����lդ�%���f�6��� f�'L�}�4)˙���w�ٴ����Ȕn�n-Q�<M����|W���$����m,z#��&�����V��&�:��T"�+ĺWĔ�x��`v�H��J����izHO��T�VJPо���H�h:��38Z��P{+s�4�*m�RX]��`���7� D�~&�=��[��0.�h,�N�f��c���+�W�=P(�T�� �(����6S���#$�����,\��D��%h�K���\gI�x�PgV��T�Ӵ;�*��Pm��o��V��-Hg?	���Y�Ҙš�ı��w]N����������E��s���r��dF͇
����6�`5;  3��nM��ٕ�����i*]�S����oU���2�\ӿJ�oq���p)���*w)��'��z|#^lvio�:��i�}c�H�d ����9��x(;`fj#[MF0o<yv��b��~��?q%P�/�Ytߛ��/�����.�|���_�*M�Ű���$
�C�`����C;���
��H�y`�3�h�x��%�����c`�T=�,� �DT�8�71�G�s�dZ*�%/	E��
�۾ o8����	�L0'����J���vY6RPG�.���Y=4O1�3#q������/x�Y$�|*1d��/�#���>���~8dC:�	_'�}�~����lP��> ��^��{�2�?�L��&�n[���^��Ա:����z�#W$�6d�)�iM��j�Qsv�!���ܩ0�d�����;n�L�n��Z�Nk��{L�[Q�bRd�rx,*�OZ��Qq�����<M�����.Q6�6H���R�`�?�6o�� p�E"��.�/� *�8%���R R�M��!���TϬy�h�X���tI���4׉����&ΥT��(�ӡ3+¤&����4��s��_�8�4�"?�!��E���q��t(1{#n&=n���/J�MO�%�g���YH�cTQǫ�� چk��UJ>Z��
os6�2�}(��]�ip���b�rX���[��+v���ږ_k��+ ��v�v��|`o>-�o�H��z%�Թ=���S:֫�&��P�UЉ[��j�i�A�����v�ſh���vZZ<�b��Њ�O7�D����o�.b���. ���L��09�}�t��,`�(��B�6Y�۵o��i��@7*��э|���\���;�w��Acث�K� j.�K����c�Yj���	�x}��
� ����q���ۼ����ݻY�DH~�#e�� s_��3�Y���"'_�D�|�b�r5�,�lS�8+dD)]�RH�E��'�ϒ%�E/�%b�9l��������K಩ [�{�-:r�^ep9�%�	�a���X���q!���d�t��ݸ�\�Ti�w\m6�|J��5��������DW�<�V���Äm!c��k`� I��F;<��)	u$��<�1vw$[��!l9v����ݐ �C�P��Z3{��PtCޞZ�}��A�\�:�*���"��u.�j�����݅}�V�lcN]Ƙ�������4�M�������i�:���o�k�}u �濻���%ԌO�M7����}���M�ʂAl�	^�=h8Ę̈́�N�@x�z��k���'���T����o�acl���C�*XXޒ��z��"ȸs���S)��I_�����*�����%����3x���-V�2r[���G�(鑟/��v��=8A� ,>�}�J ]h��6�#3	�u퍓�El�7��p}]ZY�.�S S~1���iy��`:�H�o㍇��3�ݳ����R� Żd=y�?G�E����<��v�ˏ�R` �>=�
���*�������o8���(
��c�a-�� ����b�8[8|Q��o��AV�k��o����"<a��l��RSƔs�a�`�l"(E�^��CgR��|�B����Q�H���s\!���,t��}l`^!���,��j��fDE1o�,-(����e��煹Oڴ C�JM�TJH��W1:aL�I�A��H�Q�Jך�j�ӪH�h"��u�I�=���]��f+͐%��)8ֶ������@=�-��j2wڞ�^*�L:�����b-��x��ߌ,��mZ��z�E8��� ?�&����w��1�� m� �V�T��	T�#���%_>�.��Me0Aj� � Iq ��q�Si���֏����5��{W(��U�`D��xE;�z�i j�x��툍�1r m5�~-������x��~+�V�V��Ɏ���vH��xEE��7���&�F��4�ԇ	z��2�-�a_	�Z�e�=o���`�oD?�W��?s8	e�m:����� 4]V�%'�^T�5'F�A�}p��|h�2���X\E��ЖS$�P�������uN���k寥\�9���!Ȏ9���

]���́��?Su��Ԣ(�C���̦Az�:�ڽTCU)�Y-��w��HͬHBQ�X;~� %�~'�fČ��YJd�\�����K�xi���cY�i���kD��U�
L�:�ȗ�O��U6u�u���������4~uX5�1�״#
�� DOD�衱��<5ue��X��gX�!�����%8[Bۯp=)2���4u���$�\�+^}+fo񣒃�=��uu����H�HB�$*�j%�N����W�>�O�_k)j�u+\2F�(�ϧ�A6*z�� �?�1�kc��""���z��yrZ�Y���^��� �#�j�-�՞��[�4�]����v*���w\�8`Y��)xL�[�3©�z�����{���%4�qs23S\ͯb-Y���V� �\���Q��0	��0�5��,� �[�	6O��_m;Q>���`^#A�8w�)������nFy��/��,��2td:�^ϡ	LT�+����"f�(�X���&|p�]�p��<�G�x�$3�,c��5a�D�{='�P�tBa��߆Rj� �yܢ�_�R#��]p���B�/�c�z�{0�� `1���Q��|`�����x�X���#)F�3!u�~�
�O�5W�jB�u�����IR�K4�{.��/� >^OF[��X�0�b��g�H�Cޯ[��3� ���l/,Eσ%%�J�����%�k���k��� ���Y;�Ț�E���3�S�0�DG]��,���bg�K1B�<HhYv�^��JB.�y$x]�w��DV�^�\rMKzA��K�~���T^v:@��g���QiQ�a�햙O�<�	<'���)��Z�c�U�n��S!���90G�X8�
�@:a͋d﮽�
z}* aL�nJ�� %� ���6���k���
�w�l�
������)���Y�h�AX�k"�~�$��L|���E�G�5b5�y%�"ט^�Y1NDد�?�n
@g���.�7�	g_PLm��|������j�%��9c*C�k��c��������)oOPInN$6���c�M���chzS��Y�+&��6���vF��B��c%��'�����3��Kzy��*₇�@��A�օ|�ugn0#b�H��mX��PVql/�+{�$h�rKy�S������Ǝ����hh��yB?`��eU��c]#��į�CI��/ŕ.3���}f�������_���h�,�sP������xj��:H	��"�#��O`��H��}��e��<� �-�"1�n�yV�4b�,��v�A�+�!���+�Է|:���`��6�"��nzp�^����3
���<����,���ѿ�L^#;q�qT"z?����Ͼ��oߔ���gV���F$��I��99 ��Y~�����r�AZ�l���x1^��9�o���$�% $Q�����xW̻:o0��UyKpQs��/��	�5-�����͟�z蓀}X�O�ʭR��y���ğJ��`��6��)��*YI�	x��wRq���b�����E��'�2B�r��A�]aU9��䂹�行�&�՛g�8E�~�Q7/j �pm1�l���]�k�A��.����
�*0ʍ��90�]�0�ǘ�0��؎N7����\0x'<�?���P*Ӧ�+t����Sf��I�~��칒J<x5#����{���).*z��.�������N�+�7"��!lr�
<N|g6��ݵc�������ǫ��'��p�����\	��jwQ��O�KDݧ��+�� �D"�;���������L���#��#�4?+�w�ư+\<b�TH�Qj���VjV�L�"R����^O5����1�Ϙޯ���Ud����,X��d����T*�
Z�\���B�{k�ހ�e��e�#T\K/nږ�ӳ:p��WI0�L�Y��1����J6��F\���?�D�܈�>�⃟OY�3HeI�)F\�=-������(��Sf��u���y����$�vc�GHr������mf���|����Q �{vǰ`���.u��bЀ�����j�n�����VR�c�
����IIU��g)}\�[�.��O�-%P�S�#�*7趇��*�}?���>�8�'ݨ:���,2ȇtɉ��6D���c�WD�t�Hw�y�}�� m��E�)�d}�%󬘺�)�a*�l�e��eh�փ.Jǂ��@�\�7��Yw_ÝQ_�%
�z�S8�w��6-���hz��P���X~y��\�u�jᏵ��&��zDp�S,�GZc��F;��v�D�@� $y�QE"�n���u�Ng^4�ѝ��H��kT��h�q(�$�+�)�G%Zzr�Xƈ��P�/-F<`���[�����Zm�
�,����è�S�?[o�t��$g{���w�[�B��V_�6��
���#���n��W��:��>2�Z���k�֛Uo<¦੼��M��I����A��0�O`��S�����R1�#� ����D���L�}V�h�	&iK�>Ʀ�p�Z:��͒���x7J~(�C�<oX�~U1��sӱt��.�2���y�� ���hdz����Uu����+�ݘ�C���Q�I#�ʭ����]�w�l�Vjh��m)KC����!�T�.�I�o#���iz���i����ˏ{0D@��ޯ}�s$mUcY�m	i�I`�R�j�H�X�0�nE 4г�q[�������:�x����X����엧�ͧt���P��Z�T$�Xj.{�7�Cyc�F��fV&)�ľ��@��E��q�bm��)�Q�҈#�x�m��r������v��m��·\5�Q�=�c�T&�������r۲o
��p@um��g=��9�\��C��qt��������
�+i�/�h�����z�&����5U>�t��G��f������y�ت}��v2@]u���q�6>���r�%͉JH�|�Vή9̈́���E��d�3�EԜ��bX���Tv8/�&�F�O�ڧu2�f�pO���'�G�)�B��M`3E^�;�)I���[���q�a�he���{��'�1+<a�p������(�߳���hK1�C�[�Ą�N6 r���r*H9���qg�Pp�d�(ZD�Z��f��_"��np�y����sr^B�B�$} 3k׻��-Aĸ��;g������	�R��ҕ}�"�8���fyI���ɨ[�Y����)r��q��Qw`L^��ܭ�:\,�sw>�hyJ��(�m����	E+ˢɵ�S�Ci��L͹��0[{xcD�Z��Z@�}��!�d�����f���M���W�D�����Ǭ�;��o�<���K�94��pj�����k���տ�`���?���D6>/������>�j��H!�bh�>���lS2��j�o�RT�pb��V�>�_A�0���('_��r�����7�ty*�v:�o2�W��k���9�.9�>���28��s�~�����M�ka�hXYGMa�n��.舉�PW)@F5��r,�[aA�k_qF�nAHw,�~HIBY(�E?P5H.zoвuz�M����s z�����ޯ�E-�1,3;��`	㎟{gnk|L��� 0�\uSK�ڸ�����¿K���̽�B��d�a��$�(���������#��*�!=� �s2K+3��ɝY&�]��fWSK���|��>���_��Ÿt�| �����QJP�K��s��^��5���q��&4ٳg��ծ��ᖣ�Vc�y^U!��ԝ;Ѳ�� y�PL�CR:L������r �Yo��kA)�^í4�߭�3c���z�U�K��$M�(�0�E2��0[�o�ІP!�2�j�~�\�� �T-���Ǝ@�'����#ۏ�=2���f�"TdD�+��G��4m_���}v�u�pV��j.���U-����"�p��l(��'70�?72�s��R���C��`�Jھ>$�>'��yĥ�HknW�|�X!.BV��T�=��U�[hx,a�����^����Q}bj��Y_����1W0�+�a�#�ś��i��P9��+����?�P����Wׇ���:s�����Ό6�T�r��n�h�bh1Y
�K��(�rd�ji+i��ּ���m Uf�!�	~�y��[�@�/����h�^�����16B2π�@_�V����Jz7f-���+�#��p`�Q�����S%:;��(�պq���V��|I��T�}=[�N�P�W�Q�&�����@��_���WJ�70U����W1r2<�Pd��4OfX�m�e��Q�� F�}p��� s�k�$8���lC2��(=��	Cݮ
�=
�b��e�>�
nGƼ��8J��L���f&��Z>������)�g&���04Q;Iq�������+��SL��R2����9j9���Ӟ(B����{[���(�5�@bF�m�.��y�{M�}�,� ��_�ʯ?��:�)|}�_��6���9Q�R��8쉀xI��Yd�i�5� ����W�U��c0�锷!���er�ޔ��(a)P�2S�krh�_r)b�HjN� ������+������5�*�`�ާ����h�����(��Up�iA�nA�E��9	�^��3#�E;�������v9*>���DF��z�cҾ$Vl���0�F��E/}�B���>�w�?"����ET�3!`�.j���J�Ә�]�\
��^���3k�����%W�O�
Mې�o⶘ԈLp���ܴ[7x~�N�˅'oHƯdk��^θ�+��3�)|���759�&؟@��"�ֽ�o>��L7�O��ą�m˘�`T��5UX���w��\��J1e�����첲�o�3�i�K�+k�q����a�{tǿn�ډ)i�5��b7�Y����Ŷ��k�Z�ev�sJj�m�D4�cB�
479āH�� �>�ҕ6A��/�>)��~-Uȉ|j��P�����O�]��P=2Η��]��=ϑ�m8U;dW�Ҽݳ�}k��b�@����Ic?^�����]bO8J�5 �+'���#����[t���oqk�Ύ��E�A�`���@,=%�K[��Lˑ'^i�{�iPi v��fO�s�c8��<Z�Mϙ�}H����1H�>H��|)��
=�rJ����Bm�� ���M����B��Q)hdc�o��U�D=7��ny<{{`k
�9�L�@�e:a6���h�埶���'��1�	G����b�u5�^�l\���̊�"�Y��64����f�����Ay�ThJ�,"%���^���8m�Ӕ�O�Q�K(3��Z�p�CG?E0���� w��o4O���}�&�qw5Y4�;�K��wXLX
!�>�`�s�ՙm����:��.�<	��U�� 7�f-���ܙ�SB��+R˱�H��3�٧%�>�z0�A����^�3(Iz���DBW��dY"�|VWW�6��p�3�J�nz����+N���t��7K9�6�]��)68�N��g�"�	қ��«u\<ye����Uu�=�P���g�I)Z�%Lf�X*�\>���>�}[�8�'���ZT���܄�,j������)*���j����4z%�n�aǚ�qje����Ru�{�8��w#[L�Kl�Hƹ�!"Ձ��9�/�៵������!b�t��]a���J�vZ��~�{o�Hϳs�F^r�pb�Ҥ����1>���KIT%9
�d�A�
\�@����������!n�*-*�U����rI�}տ~H̝�ZB��p�#B9�W�Ƶ�7�����2�`8&�U�؇l��80����|�/8��_�H�E�EdQÚ8	�c�\%FC�[I�X�0������w�eF;Cg���څU�-��r�
n:�M�V�`�t�KE���R�CΑ�~!�?O2f-�=s���S��$&����8��"m����OaiE���Y�g�иIq���NQ1�M��z�݊'���H�}%m*���:`cԪʴ-46�����:Y�N\����r�DCShO�X��w�[����'f4+�sn�P$���
�h ;a�<�������y[G�P����)�Ei�� ̿`W�a�Jo�����0Z��G)�$��|��\Cύ^�z��¿Ac�[�HFZ��߳\�/L������$��`�i�����h�n�� 3�1�N>��u���<�����yb
	��h�G83G���	�àǍ(��|v��b�t��ɧ�3�ճ,&9tq�s�^Mzt�b�|	��[ľ�;[�)�ѥ�t��&��z3t�K�����ti���i��t�ח�6Y�!'끂�1er�?cCx����� �Fj���2Hu���>o!6q<���&`�"Yҟɥ�ڷ�A�D3mnTY�g� 
.tf�Y\�������Wn� w}�I�Jj��J~���)���ƀ#�w�9�9��p��qe�p��u멊����Y�
�#i�ǫ٧U�-�^냎�f/&�#���/1*�`���LSس1�d�tq݌�K��8f���m@�(.uL��V|��'���T��њJd�m��SK�/�t�[t� '�a�m�Ϸ�+���Q������~�}�MF,f��i%Ni( �,q=��=˸Y�fc@2�]�m�y��V��(�\�U��3čEvk�W�f#'&��'�(nx�U|������@�K3��Ӛ,�`kJ��a������g�3��Ԝ`�!U��_7fꬆ�����J�!����y�[��u<.؅Z������Ä�Q4�t�����"�7lw�JhL �
:ܝ>���q%���v�(R�k.C�^T옼��Q��H���j�c?��2 �:>I��n)Vk�^�:�kkx3\�g�w��f����}!]e��φ��9OQ�t[t�*�63�L�B��x��4�ɞ,���`(if�FX:�}� �m|���meΩ<���}��N+nn2�o0N���N�n�j)�w�>�s��^�sm�#��H��[׌~]��J	E�\��Hx��c�7a�m1Sp`tş{?!���JR��+*!��AJ�]�]ĠF\��T�|�di���)��mm�RC%���K��(��2U��ʴ���]�U(J��4k�-VE�<ګR�ɝ�?b�^;û����[����$�p�H����>X����(�T�C��*�� 	b[6'�l`K�~C�V�Z��tE{�$$ܽ6xs�i3ٟ?g����Tz	eIy�"@��l���;�N��ꈣ嘥���e���FWV�����"#qv��:P�f(c�GT�<v���Ew��S��%k���ɿ���ܸ�D���TD������4���������gR���:-��Cq�޽�h	k��ʮ�zQ PRq�]������|u�Ż��ARXEм�����L���ee���±L��k��1n��cQ��Rih}��ú�ʲ���<�[G��}x�M5�d�:��L�Dy ´�O��/�r�Z�F��Sz6�n�(Rb�;̧E�@����U�.�Q�a{4�|�d�H*�J�t�	�3����S4��t�z����hw����e<8����S��������v8F���`��o������U�k@X�Y���ߐ��Z�N��U|Ǳ Qo�`����6���

?!ؗBŗ�3;P����?0��׫�!ʃ9���O�~�4@� �$>��'��@�\�ȋ���~��[�B7���e6�����Ӳ]�����zi�E��2.iEg�)�ҝ�GR�ޮ�a���E�CG$���.���tR>3:x���:����tP">��ۈn��>͢
�ت�i�~����{�-=��3�E����%���)V@Gq�D�����Ч&�vl�|.�b�ौ�LW+�b	<����?�!������j�HHiC����b�'�����22$�K7b�k˃��G���<��^B�
�w������J���δG��h���y�[���mC����"Z����'=Eg�*L�Z�=@��-�0�ܘ�'o�L�:wR��]���nK[�խ�C������=Ujzӟ[h����O�XF��8�e�e�RE�?��@+ _�G
���G�2�S(�����;��r�}�C��wܔ�ҟ<����4ﻸD��o�e�����i��hq�<:�7S[�j]�G4j>.��p_+�*5�����9���[�+H�W�bW�|�9(��g�C����*����<���7�>�h_�{�GR�m[�G��J��uM�k��	�	�Er��1 T�q��*�{LY3���$�j|�}j�UsJ%��T��"l�;B�/ܕ��#*56��`'Z��l��� OvG�C�Xj����{Q�353l���cS�{Qt��YU�PGBg3h��nk�>^\kN'5�u�9�؍f�o��5_1B
d���
�Z�4ũ�
���={����_���3������iO�<�^}��s%g2������z��Ω�nõ�Z�'����4I���44Vc����b����m���E�4酄�*�|OsI��ciG��N�a��i@0�yP��MyI�h�`�e���:C�c�Y� �K*��z�p~�{��Xm@՝l��˽mq'r�_1v�N����~��7�)N�7�~���/O	�*h�^]�/��rv@3;q��(��b���X��k�v!��+C�My?���lo��������M�O6�aʀJ�ا��u
V�K2����22��l)���>GcL��B}�8z�P��b:Ae�5����7��+�����e��m�F����$l�S*�X���v���Ԑ�KEs�`�x$���i-��� ;!��CԦ�fO�T��i�����QM�?y�,�8�J�?�K�$_��E2Y7���fS� �|�T:��kB	��[�k��[H@:��P/0� �u���Wc�"����%~w2"	�#}�Ⱦ�w��.p�����4o�J�p��$�B����i�Z��8�j��H�n~=���Z�訟r�KÍA�d�|Pv�^�"��:�
|�C|�-_n��G��C�*�`#��_�j,��WV]L3
���h��/Ӫ�'枳o����Ͷތ*Y�y�����N�p��@c8��^������mB�9|d`g�����U�`NB��Ze|%��H�0��|Ó��i1/��p�6 ߳���b/*�Oc�6��#�E��Ҝ��e`l��� ��C��t-����a��ƚ��C(l�a�g�&����107k&�I���5Ϻ�(2���F>�A-_���W�:`�`�7���a.�YYēG֫5'5�?�T�Ͼ>�lx4�m{�?����K�gC�f�4]e�z�X`�}�m�E�PWfw�NϹ�|Z�GAȬ��.�u��p~�
�(�o*2 �U��'0���,D��|��Z��!�L������J#ּ*�]��	Дo	��5���F
��J����
j�W��ԟn�K����QF[}A'O ]�C���q���2�{�;@QG�gu��M���|3�-��*��*ii&gf��pC
��.�L̘%&!�>��L�r���&�o���ū�4��H;�->mZ%��]����y�7-w�����O�����8�:m:L�F�I�Pb�R�C{?B�������'A���V�F����vx���_��$�?�\8|zt��4!���H���t�g�1�W8)!AW��*�F�x\�'YR�9>��,�"-�r��,�)�j
��� �����@D7���Ov{zx��8���s=Ө��D�ԯǰ��Ƒ��W�b����(��)�8�K���q�I�)��4O��.��üzU�I�>H�nq
Q����%��Yb�;%���(t҇q�@�ea?�B@�P��4B��V�Pp3ov"�fv�L_dv0g��W{��^�%c+���_�B�׋�=(�ȍ�<�Zb��ze�1�� ���&���P̧���泮�$��G�9ȶ���ׁ���?̚��e�i��o��ٓ�?G��+�I��n�$�Qg����&��#�7�Wϛ�۽��sc�K[! �믾��5���sA��G%��k�b
�m%O��,bU����3\�v�ݠ�¸�)j��F:~�𠃷���0���tM}�x��J���v��苊r��+$>� ����"�x��k;	�;q��qo��3:��&�KP���s�z��i"$�y,�;�v �뀮��l��	I ���w�	����Y�L�-ȏy���sS�Mҭq�I����+E��q%�gi�C��>~l�����E7=���D1���ɛߔ���F��c��jE�Ozl���f��`�3u3iX�W��fKPZ��	B����qE����{C�%�Q��rr�|�O5)����_�icj�ˑ,�{B�������ڼ_���R$Z4�U��N�TP���LV�8����zF$A��$�*�Q��	;�AS�����!�w�"G�ҲF��:�T�����4���d�2�t��DHD���� >ʐ6閛�PF!��U�{Se�ܞ׉�C�bBm�3PT��-�8W5�?*�� �����|�,�Şs(�G���.�밻b��n�F]�|�q&�zzK7�*�G~�޼a3����E�Q5��v�y��RՄt�����䫽%Ѵ�AzW���,gհ]�-�t:Q���e�zi[5+A����6J�/�
���Zm \Nl��4+Y����,kY���V�<�Cl���sP�%v��A�2F��i	?��l3 ��b�X�S�:T��� �7����õ�>�����r�fqZ�D��N9��|�J}HßG�&:?j���HK���r 9E��X�^Y�*�{K>��붳�f�������Aބ��Η�M���H�Ĥ�} �L��ҫ]ɬ�ދ��5|o�'$��B(�D�*,������J���WOP(2�J������w�y��m^/S��O[�&fB=k�O�֍|��Ya��^l���7=0Ĳ�#��f�Q60L	&=�� �9�7��������7/}G��G?�붬]��U�;pH2�oz�8�)��
ʴ�-�����@��.	u�Zf����ɀ�&H�;���-n�l+H�c�b�^���4 XF��,������T(��� �O�f��̶�#8*a)x��ϗ������7�z( 2n1Q�s�=j�Bv׀ȺI-F�&�BKU̝C����82�E�����hQ�"�t!���F3���	1e�{��/N1� �A�}n7��w���61���ܴ�ܙ��Pk���-2��k�?E<ﾡ>^��vb�f�0�ͳ���$�Ks^����X�~�A?V]���~�t����"�;e����U��=EW%x��}O�+��݁�8���8O]�9��u'F��2qO�wۯ�FAG�*w��tcd�y d�2�L�3��n>�虳� 
 �Kj��\dZV?qX|<;��^�}����GG�;�%y�y��r ����*+Mx�S�&o���CW��M�9�w~H�*�<{ܹ�&\��%U	.ߗ���ܔ�����!)9o̠YO {h���ۣ��B�M`�2�>�+�����j ".l:��N����kh�>c�+SV�lds�[R���������:�l=��*�)W�@�ju�{��������o���B�}�d��stJ�����&à��k�ѱT�::��6� ܋A����`���i ��2 $Ѷ:�Z�}bЭi��A�T9	͞�6�Q�m�<`)��[;A��49�k�>��q�:�n9�4\zQ,u��!�*�h+=/r������OHn��)��-�JΘ�7�\��a�P&��$躼جY �r����[ǀT�>AVJ��T)�
�M~4+J�i���aP7J�i�{H�[��ݷ���Ag��S�Fy@o`��Ю�狰�W�X	���E����r�%�y*6�AD5�L��W.��~C�-T�楢���$� ��✧���q���P��]+1M���&I�'2F�@�A��?sz��@�&W+�wR���̃�.O��q[ AQ����ޣf5�c�Xm�h��;��P��*aO�?��˟RH�oj���;����ə]�A7V�a��Os�lS5��PT2�W��.�Q�KsQ+RqC�DR�[����K{�� d�E�h����A�c4���ˉ>�y�N��(t�/B�	�{G�MH� ���!��ދ`3�	����3>Q7г����TT�v������,n	5����P��w�-��ZͅF̩ΑK�s��~�!G���d<���aB7�i�޻4�Gn�����aVYQ��/�j��1o%#R+��C��m�uA�|��=�>�8�mZ\�J�i�c�N6u.#�@Gw{������)N\��D=�GMD����O�JzyhLEc_c[ۗ�*ԣ7��/N���U���s��M�-V�X��Y�j���y�/�X{wa5W�w�p�֮��.
��~8Q�#V:���;dт�b�t@������(��z*z�7ɂx�Ѯ\t>)��7�Y���tcBYL��ۑ�6M�7%)�zG�V��Ћ9r��2R���pMrFlW{�5z;�t�ϧj�]9'R��!.����ocժY%m���+���P$��o�w���4NG��	�|�J�}��drѩ6F:��3�(6�,�0��gg�x{6u������Lm���4��r]��u=`e]����e䋴z�[�͎-����SBʲ��)����8OFQٺ�q1��H�A�;q���j$��࿩f9�����l=<э����,m-rk��HӖ�O���{1K�M�l�*䞰�����s�/�	�A<f��"�2�����4�%8yA�� �5�ῆ3=T��q����ZQ�?�p^֘O����:t�W�eȩ~z/����gjJ��z̑2]�%TY�ʲ�r���K�8&��X0SO�����ƹ�8]<:��t��ɂ�x��@�򓘘E��O#���>h�?emR�H�{)�H,�ɖ�n���5�̐"���� J_ ��y���W �W� ����\��F�Ǎ�0���f���_يi5�EXi�*q�������0��}����e� ��5~����}�)7�Ӟ	��F��%5H2�H�F�5�Fl<m3�`��8;n��҃��8
u��h���la:���u��4]q�4={��[�?O�ɚ��L5�-dB�G�Y�M'�G�Sf�X+.����0f��'�j��|C��>F�=J�.��eԓ"�K�YǦ/ÔIO��,�@����iE�'�R�%� ��@�`�^e7������Ҽ��P��#7�r�����tL����������?"����f�v�sTP�mS�Pq���Qw������,��JR~���^ÑxN�bI0z[��s����bJ��m�=�����N�d�]�]����o	^�m�BHU6�A�-��x`V���ޕ}A�i�ɻ{��8� {�v�1[ܗ�+)�Vj��f'G�
" C���}h1٭��� ���:�^����d���)48ϧ��K�&=ZXm��Yp��h_;�;��K�T�l��G��ѻ�-Q#�M� �cïtƵ�����8��pu	�?��PE������a��]�j2Q��.Y��r����n��m����8�x���W]��ع����ou�|�{�j���u+�6�UKyb�j�>��Z���/."K�O��U��P�DB���Na��	to�P��Z(���4�4HP5{P�fc* ?�i������DL���f���U6u��ƽ���G0���eL�2�.ir�X@6����+�4c�~F^%��q����CJRibe��ozA�� E�Ư�v�U������	�E)���	�Q�E��[	 x��F��|E���d�K�%��p>Fӑ0�E�=ί
�;��j��$cI@v�/E`o��I>���·�`��٧����p8��LM���N��v�b���y�=�:������ ���	U}���(�/x#��π��d�O�Z�Se%��}��$�6d�Z�g����M *��r80B9�;"Ĵ�ó��(��4���6a���ݒ�8��雃<ǭ����v���q���F�lc]ov�������[�|�!ؙ��Y��Y1��hM��;!��%�����(.OG�����Fb	��ݤ:j� �]V�!oo��I@�>%u �C#r�i�	Y>�vy��$���99Oڑ��}L�Kln�7�&��I ?ҷ���o�@�����|���y	�H��[t%��h
	x�o��j���j��(l�M�$�q��w<y�����C1^2}y��;��ӭl\����1���wM��x���Y��4�4T�+�uY����%��`;�#�%<8탢t�4
�������^N7�{;�ѾH#/�S�yl1�'���2�F�V���h�b��`��ey�}$��t����R��LF�n�gp� ����=2�9�~Ŷ�Cisu�h�i�$�\�x���iݝ7��r�c�q������q��U
��W��l0�o��Fg|�=�˂�d�֕�ߓ�8��y1��3�����m8���y�gq�0��Ev�/F��'")tM���*'���]�+�)��6���O�T�]~����鋗^*�7m��V�b�'&��(�*�tc�(��Y����I;��AX�n�-\�}�}g6�ߥ����/��.��]�/�� O`.g�;E�o�"��`�|g#'5�͗�>�y�u�Y�`}ש	���0V]�8;�ęl�B}��_�*Qؕ�y�<���6���w���˵h/%L�����a���X��l�ps���8�!)ӧs����Z�pe�ߵ���ik���k1�s���.p�w�i�-�~廒u	5�����7��A�?^�qM�N,��t������?��m@�`��Aq��P�(�DAG����\��[nʈq��(�"���#cLa����MTId��/&K��?Q���Sw��v~v��h�D�I��9��-x��ѭ�_i���ِ,��'v!t�=Z��l�ťL�F +�K��K$9ȿ[eO�q��K��<	��8�s.Oŕ��uV��d�����"��=�?N�}����&K����񨤮�`5���
l��n�"H��M��xs6b�}r����#ʿݗȗd����7IX��x�N���{f�Ą�Q���^"y]�u�
�A�r8�׭[}���b���z���C5�( ˨����^+@�ggo�}�#JE��Ƶ�D���s�Cj�>�xB/����e�ؼ�F|}y�f7����X����ԱZn���<>��I��3�8b��VkWu�>(�Ӱy��?ܑ�z�\�����<g��uX��g7�ROes��	K�_Ǫ�$�a�����Q��ǈ֘����j^P��#p���P4m���E�C��Z��`}>Һ��W>��d35(l�M=�S��d���`����rhb���lG�Bap%�"m� �����kC���4��2>�C�<�׊x�����[���AY=��	g��@�S=�7{�?������慡
;��j�V�o�0���3%t���5����~ʛ��=�)$�ٖ�	lЮ/��Z��h/�1p��3H��y?����A�%5����;
��N4����0�����!��rk�Z�Io_U�~���sc�� 6��o k)@5�:io�+� _�X�hX=P��e��Z5.�ʯ��Z�w6��Y����l�?&���i�(��u���^�Y۟g�).y�MHwv�lK�7����aؗds�!Z�Y�� {ɳ+��}��s˘�3B�	h���`"WX�V4i�Ր���>�*e�S���P��Y��
Y-:pn���&�G��4	���0�9C�K�ݩK� fE�qq��u��4�A�kȌH}�bj��t�Ь�9���׎L���-`hwM޻H]�z��hF�*�����̜f���.o)~��C	tLc��"��OJ�Y0�DP�IQ.�RS!�+ͷE���V:���)d)��oVOB/Eou��t<K��Yd8?�̴��l�
�%�.5�}��"�Rd2�n���ݜ��t�mV��f%����bE6������5 (�r�p����Dk+�$��Akɝ���{d�M��%���C �P̪(�u�Ц��W�@���dl\-�D
l�1��è� �#��>���sdr(L�&�(��4���Q���7�^��B�������U3�l��=������Si�pX�4q _4�l5�܃�{1��w�q�O��n���T[w�L�O� X;7�/J���y�?r>!4�,��N�O��<�%Z�TIK{���7���&܎����46���T,p���)�{� �N�q��/�ɽ�.'\G+H
I�Ӣ��d^3Ƹ�mU'<i_��m�9����\��Z�Þ�ha��N=�+ ]�)�r�������v��*a�0�4)/�/i�3���z�[�M���ݔ��!�%�D�ҕuG�� �7^$��\y�c3yh�;�g �)���PDq�!y}��d�:
r50��/�M3R��-�'�+�X�n�'gd )m|�W9�A�|��>�.��՗x�D����D��R�#�Ny�)WK�/fL/��y��<��!���y��=�Q���m�?�}�������"{w����Ϥ�_<��-x���+�Vd5�	`���	�����f�*n#ؔ�d��!_�Q�	�V��3���<6��?��Mؐ:���Y����RQ,���C5��g��?���?�)����������D���S��i�n(��p�A2�N�H���g��6���G9��R��EH�S[����Yl�&.V�&��qCqa�ce��G4�	�o����\* ���|(�xCi�[~���"��Y��n�[��W+��"��ȵ h��Mx�g~j��
�Քx	�a��$)�eRy�2O�12���	~!OY~H�'��T�9JY�o�o6@�?_��KֆB�Bd%J�o~�6s�^XѺIm��l�� (c��m�B��9�Eר��E�-8��Q1�07>A��(�s��Pd9�jv$$6I�$�ćZ<<q�C8w��[�S�R���{�L�,Zr$x��:Ο-��>��鍆0�P����j�W�Qgi�@Ft�.�����eY�4!�.]4k��PVII�~���$�κYz/�U�RO��6�������� ک����p{����ZZ&XPW{�x�i>�W��(`���Cb���O_����� �X��En3&VT�����H�Eyq�~Z/��.���.�7/�S]�B�������~��@�Ӗev��E%z�*�ͤ6.o�T��v/���9&[<n�����s���P7>��`��A��kl��gNPY��/� �<͜��D�K7h�G�*$�nw����� ��]��tνT�h��)��ɱm�OR��|��^y��W��v�E�`��J���<\�~�s��+ޮ=w���R� �ѡW{Pwj�T���{�D,X>�㬠��![}�� �Wg%6�����OY�"";������mB&��56f$''+X^)w��4�ƙ�Il{���S~qk�2a�S��w�Ƕϊ3��1R�G��5���7ʆwN�|Y�+`N�8��ϯ�+�ݾ�=���+��ᕯ�r�O[�UY�sOal�c �L`�ڧkt^--� ����t�c���^�n_�ݜ;9w�,�昀�t<e��̀K'��`�`�3tE �5W���z�N暒ag�MA�'��<0SoyIg�N�M8r�A�u�G��������U��/��mJ���&�?�:5}��	��&:yyu�$9ޢU�-���.��� ���q3L8b}�Ơ���5��/K�e����A�z��yb���u
�'c�p8��{wt�2��{���^М���ʿ���Eu�z��Ev� t�t��u5���Ω�K�q�bT@������mZ͢�!�Y��<%���%C֡@��d6Yܜ�� ź�<,[+^�G�Eߜ	���9� B<{��&�ű����4��R
NS��ة^�>,ry���(q��w}��լo��hݩ���'���\���{��,�l�9Gw�|P�0@Lx����/BH���oH(��L�6y/�{0g*SE�rVsm?جp-B��l,�CJ��Tձ/z�{b�߮a��+����9r�R��'5�"O�ǟNUlJ5�|5?,&G�4���
��ٸ;�>�ϔEH��̛^�÷�?�x�-�e9�!�=�-\�|�����3hP��D�h��6FȨ�zeTUȩ�9��*'�f�bT�vzt�Ѿ�"7L%y(S����e�ѹ� TH�вV�/��Y� ��5.g��uO��0t:}y�.l໣�O�����9b`k�99�̠�?(�M$��Qi�u��$��$+�s��,X2Gp�:X�C����m�P2P�g=zj�A�l�7r;(�%P��(��]��	V�� ��\oq��<|���um�&�!��V���Y0$qv����ms,X��D8B��qƣ� �cO/2���𺭞����L -�`���7S~�k��@.�A0�Ӫ#X�ʓ/�Q��0�G!��&�=�^��d�hI,0����#�D2��j4��h9��d:a(�瀨�q$�F:�eV?	Ï!�6�W�#�]�"�{%%��� �
�@B�K��MR��.����ē��M�!~����p:��{��X)����7�ͷu�vc��?�L��rJ��B�6������4��*�j�X\�M��T_?U�({�)�Hg�x:��y�c�"n��gm\v;��vk�~�˟��1��Sr�����Ꮁ�%��i����f`�t�b=�T�$j�1_Ҟ��Ы`!q�Q%��z7����e�!�2����6=�Y�3@����y!�%�@��ѡR�k��zo�/�+`Q�uc	��Cv���ٗ�-0����j����[ʀ��fԷ�]^<E��]��\ �����ՠ"���nw|�z�0|�"�M� U���`%�7�X�q%�;x�|
���X{��[ ��|K��,r�}�I��Z |�i���ĸ)�,�؎�J�#�7�����䄤�
�|l�İ@0m�|���@�X����wz���p�m"e�Q{/P����؈�j!��'X壬\�E���Έ�5E����Q~�f@~g� ������m�� _԰|�|un���y���UB�@,�B �asv�p��)}\%=�T�-��$jc�ϐ(�Et
��DHYR&�2 ����.c-w9׃][`��=�)����D$*-K7�y��'qs��c�O_By��	�!��t��p>C	���L���T._��M8ȑ���� �e����\TL=���ܪ+����)Ɣ�B��$%܌>_�!����U2��A���ytb��Z4h��K��KD:�����K�����\Ԡ�>"�����^�*�`����vg�8��:z_�p����)�3@�tfNRS��ƒ����0XɅ!��<,���诔dS]$�'r���&�^�Z��+��in��JK<�����z�&�*�l!��0;�Dd;���kw�X^���ȸ0.M����	���2��i� i	�#���пO���x���c�C�bȕ9Ai��N�V��o�\�[@7$U=UnD�J�=:���ێ�������u��:z��b������{�B��w��]�Ps�:�j��TP8�NJ�]�O��d��n��C���Ӊ����|(�c@�J�t��d�%�A0� �0�6Aq��_���T`��'�މ��g?�c��z�`���DS�݄M]4eƳצMTao���s	�� �Y?���b7F�"�A���D���v#F��CF���rq�3��RW�͒����5tnݓ��F�Y�A@�n��˝�dʿဖ������-�0�?n��}i��`	��|15���`�V�&����H�.�_^|ri�ɂ���#�j� ޅ�
�\�k�M�#1ܪ�^��1��L+p�L�s�ѡ��+a�u��h����)(w:`�=��vIP���1s|�vA�/���r�sҍ%w)�-}���lq^9�v?Bgկ��r���}��='�o�FX�k��9�`QeTx|�*Ńr=��,O�3z�)>���o����KI�Wu5t�t)��T���V�1��'Y��{i�ٟ�dXz��rQ����aH"S�a���,>�I�S��E)���*�F/]��v�l5�i��1��N�`~�C	nl�l�5�B�Cĕ�3d,��ވz�fQ���<�|�\��m�@��n<а�M]k���m����cO������MI�7�lzVfS�C���nC
�~1�'�j�Y&G��G"rÄs�"���]BAؒ��D����:�A6l4�Q<�m����zn����!L(�$�f�.�2�y�������sV'"��ȎU��%)D|a�d����$��iiH������B1�����J8-��ZwWB9�L�-����.4�m�ଲ��^�c��K���;;�nρ#�U�ۣú6D�ι�܀�]}�ͩ ~�尞H���ɠ5<St�zoÜAn���aV�?�ޤV��(q$��_Wi#&�u��֔�Zת�AkrQ���O��J�<����k�%wЁ�&n,�[y�i�R���?���_z�W�w�l�l� ��E��y~�c�N�����Ƶ
9��ΘV:|\}� g8p��BuU��qg?� ?�����m���K׾1�bb��@ӊ�?ʉ���4fAb��*�x(h�]�j0�d��M��c�l�N(�xԹu�')3l<��=�S��6�G�p�EQ�l�l������E38���7�`��}�-ځ����<`:��LA��9}	�,�:����O
��1�X��v�zk�Xp�C���� � ��d��6V&��S��4��V\rCE��}��_P^C1-U���&���a(^n�L뺰�B���$���2k_�,�nq�3�nh^h9`+�rQi��Qp�����,���J��܀���!X?h &��� �ut	���ۖ�+^�m�H�����e%J�L�	���S�_R^�t��� '�^ǴZxԯ������IVbߪ^�#���#�YR|m����[�y�H{5���꒏
��W6'���.���y��uU�]��^*��$�I+)e�+l#�����3���ÞZ�V4�m�>W�9��z����7	�����xN���8)12�\��0�=���K��0$b~��s9�!�yt��
�#�k���Z:m�	ԙ0���P�4��h��CEu����e?��u���0)F�NjyV]�lbي��1�}�|(߮�)r?a@�/B��/7t!w�fp%��5�w�B�WK��\��{O�-N��"���U����*���E�#Ų�N���/���)������C	(Vh����$�aٸ_�y5C��%~2�����g��2=D9�sKT]8�% �ɬx+��Cc�@B�'�{e�3�>d��fX={�>m,tC� �O_"�F��to�Y�i�Tpͭ!�\ ��dұ�뺖:�ݴ�[�\��#��I��ւ����GN[T'?��Z�m�ˇ�F�ا�I�n�T�G�ʑ¯ӛN�ɂt�������y��E���aB��ɲ1s?�`���I��6�-z*+|�P��(;���;������<���8{"lb�H�/vHk~�T��T!�!�Y���䥵�o8��O�wu�W����P<u'�,�j�K{>��+�j��f�3%<r*q�4�KD��h�}<��sỴt��9�,?�l�Nw�8�7ѱ�9��u^�Jy��61�)O&�~��b��{ӊ��a��u7U�Q�~y����V����{A���G�5d��;ȩ����MAI�x�q+���6�Z��0C��'�����&��{�����]=��AN"�@�i�J�䖮�Oѐ��Mt���o��HAŪql{Y��ŵp?� �1�|�OG��d)W�L�:���|y���,/6�C�,�����Cxߔ$�I�_���O�
?�'��^����t����f�X�5@O���(�F�W�~	P�8�m�Z'�Y�߶��'e������������zf@�X ���Cܓ)�W��9�Y�q�#�+>-C�L��T��'|6�,���H��
���T!,�����/�����ˋ����FfO:л�Xw�d�uQw	x�z�{�L�L��Ee����40*���Ɠ��ɯ���NB��q�xW)��)���%��	è0�(LO�_hcJ
�m��<q�ԧ�����)Çٗ����
�'0h���S�^�9���%%��(83��#�Խ�ts���{�7�JK�o�>�̶����0���)��>�uU�iE��J4U�#Y�D���njS�cl��-P���v"�)�m,R���}�#CX,��գ��� �o����?�6 +����&Wi�|�	ظ�����OM�^��;�f�^t�Lz�6u�8j����np���b��8K�Z&Ɋ�Q.�qE@����ܼbZ$?��9�QV���J��t�A���٦�V���z����h��z�����p�d��/�r9b��c��n���!�]���e�سt9nT��-�U�ڊ���C���eJo*��^.�����y7D?�f�D�p��v<��b	��;�Wx q;��SW�N�����l��ŜZ����R�p�+�vj��+ޢ<u���7��< ��;�Z�Ԅ�ئ"Q�w�����v�A� �r��ͣ�����ǰ����~�wl��>ы<�V��cl���'N�K��7�hb������Q/b":|c�V\�9�6�mԇ�H&����}��v����*��V��]����J�,�V�trnGJ���p=�!���ǵ���1�!.����f #E�c+��d.6pC�%Y-I�~�����V��
b�M�(7����ſrr7{Z }��R╎��2sfH0s����L��1�4u���)<K�ҵ��OtO:����i�G��u����G.�r1�@��k�=�E�Yb������+�Dy?>{�$��}���	��?���P�S܂>��;�^yW6���b���p(�m)�=l�gJ��i�iG��
7O�H��+�k]�n91��T�]����&�#���w�S��_E�C4w��:��K��!�`]טR��mt�Ԕ��M�G��A$W���9rj$�p��cWfQ6�N<� :G���j6��p��� �Q��̞k��b#Ƌ=�$�#
��gH9+M��'݅�b+V���E��m�~ ���v�79DAH`����j_M����k?��L�pR�ݔH����ό�}�Hk�`�u��OW�㽦En|�N�.���~�q���3b�G]���y����A,"q�����Ʉ%8kU`x3��YRX6߭f��j��G!i��/s=3u��Ư,-i0��B�T�\-U���$�]��w,��2��D�ѰM�4#�4X������4�/��·\s<|4� ��^R �Dl��xt>����t��Ad�B]�`��2�-�#
�ЪFw�>�BntХ���蝍�r%e��`yy �Ω
�R_nG�F�S��������NZEln�I
 �& ���(����F�[�z���uv�R.Ѣ�$�i�Ŧ7�ȡi��^�(pY�}��\�3�"ں�U����nK��6�0b��`�aM����c�Uz&�R$>M��z�ɻ�L��&�.H�i;��Yy�BX���Zl�GD����l�ߌ,����= �G�l�_��X��xo��E��5V����m�����Dh��g�Ӌ��8����R⮠���Vx��S�G�=WTh�YҶ.��mto[F��c��ZV�[��]OHd�<b^�bn_��S���NC�3��r�V�c/-���):� ����%�6�MXϡ�	��U,�x�#\�@0ƕ���F�Х_�'���vk�]��ч�[i���k�O�1�+T[��^u�ο���d&�I��q�i�F��u۹x�.���H��O^�� ���踌���?U���DZ9:lG��zƌ4w�b����5t,�	��`�|��>\�I4�;k#ը�\J;�"������cĥ��be�ƌK"1�>���C����W�JP�@��� 3)�|�B�=������Ww)�'�3 sj����A�bb���.�Xڱc�E�bng�k�Տ��ck����P@UZ��&(��F����:�C�و���|����}u�	X�Lt�B�0�P�T�);C8����9�g�KVe�[��X���E�r��%�Ĩ��fJ/]��'�Kr��L��8�ZdU�M��J���WLd�W�ؒכ-4�F�۟���P�e�s���@���N�-��`�U�N���EQ3	��� m�CVɌ��J_�����!�֦��������4������ho���|��٫��m����1'S0���y��H���'�{'�ʳ(�L����n �ɦ2M3���uYj�5�Λ�|�X@=Nv��oဗ� (ȿ�pE�?�avV4�����%&�����K���0�)�7Жb��pHzIwGQ@�FZ� �_G<���U���Z�gi;�טv���Y#Br�-t�L&/(q)�D��lpL���}�#q��B��hi�Z�'����A���I�+݀u�Q�,�)0��̵آ���Qϧ�Tx�W��'N:ޏ��/_�b�w��C]!ʆH���,Y]����Fu�)d�:������P��Ze���GEó[HA>.3�K�[@sXj��7�I5��QƮ�,�J{e�wG��4?4dX�H!C6�������1���/�y�P�
l�D��̂�oc�)�t����y��ݕu�r�K1_a��~� Kʲ)�����B3��b"��A<P��#�ik8[$�EQ'���;A����M�"��)���#8_�+�r1N�w;���L�7��P�jB�.�.Τ��67K'r)z�?Biu^h0ЬT_��(���0����xzu�]. �~H�E�k!]�N)��  � \,�x��m��`aq�}<�gJ]O�1v��~mB���G	h��|ei�
�gK���ʵa�$��Q��[��K̾2!iG�A��g"�%$�� ����ViX�&��p�r�ܤ(�����4��:�[{��!���$����3n��<z����@0+1O<;���;�C�����{1��ܕQK�&x
��C��4�<x)ӆ�x���7n�x=���^_j���>�!@\O�.|�]nL�k�vm��7���/V�X�����$L�I���l�J���4^V���Ͷ�(`�*�\�������?`c�,�P7Z��*�O��t!�4#�-B{�>'�2K�|�2�|�6�p�wh�Nq_�[�H�l��ݗ�9�m�	��Q��X?��5I�Q�&��jߠ��&�~9��-��lb��[}\�EHl�p�t�YB+e��4���oq����w>
�����E��})>��;DN$ _�@�넒�|�����NYp{��3�*�a�(:�V��@��T��%���dY�zv�X� /x3��;�H:�ns�B�af���M��y6��el'-�H1k�\>��HR�Cd�h��P��[jb��X��=�H���0)�_��������[��m��*e�y-�3x�ҍ����GL-X8����z��S�Q9�.����I��fa��#3Aꅯ����%9�~Z�HQy��?#Nc���p3�|�2���d��jÊ�KիU���Oީ��WtB/٪=hq�'��摊AzI勃��j@X�P���F�L���G���j%sB�v��	�-����6�������H��>Φ�\�����t1.m��@o�yu��ɟ��a�M����\٪�o؈`�J̛:?8��
21 ��-�@'#�����2��ӥr�������9۹xsX�+$+���:��F��fJ�~����+�ꇓ��Ė �_SxM��X���:��>ߎ��WvΊ� �W:|-��r}%���,�F�S޸��F b�	L�@?لL�W4���e�괬6�Fɭ�����d�	8��f-��B�΃��j�iUS�aVP�z4���P؂�Y�.)Ox1W�>�_ph���N�klT^���"�~������kԥ�'�l��)�j?R#is*���a �7w[K�W��
��]��O�&�+ހH�o�������M?z�
�"�T`�D�r�s0����Q��G�2~�5@��&����u�c)׉V�K۪��.�G�4��ΠJ3��b��ؖ�+Yσ
���'��g�r�-��\.�\�`�K}𻢍m�}-y/�aU�}HB�xe& E av�� (k��VK��)Vt�|`�9Hxu������RG�����
��]z7�,� ���l��J�}�oF������z��.O�%s�{J�<BXd���d��\��O,��*iE<=�¸
��>�+��H�b��U ����1���5��,IF�	�����s����A��W�������5p��g�����m�9��Ni�`ou|�����B��ݥbS*t5l��z��jw�ԗ���ʎ�q��_la4�L�R�RH� �E��R&E��&0� �gFl�Ņ��k����x��&�N+t�<���O^<K+!e�!\@1�-���
�~^K Y��6�ݲo٣B�i㛊�eM�8�į�*ax@[,�]��r7U� +��AM�������3@���Q 1f�G�<+i����S�8"E�U��"�W�wbq�j��,�j�An��I0�m�V�d#=мH~�Γ�'��%e]�Xi2U�g5�;��I�Sl� b����p:,�s�X�\��F�5���7:�r�B-�n[/�rHbm�~��"�m��<���7��ŏ��3��c��=(�uS�i���ƩF�T�Fr��i���Uװ��ݘ�4��}�;�jv�owYc̞F�]���oT8#V� qGK v�1����@������0?�����χ]9N3�#�_du%D�w˨�97�O������3�a4�;�ﴝp��Z�	��lv 6�(W����`{�g�E&�-VX��X��G������Lf�����B�|C�g�98��ܹy/H|A�neJNY|H��,a� (���wE5rZ6�@���~�=�L�U���}k�!��9��,��c�|�l�߂��mUë_T���O�"���q�c�L���GrY���>B��0b�����{g�����Xs���E�V���nIz̵����R��?e���-9��N�x8Omk+FCQwr$}��n�+{֕b%{�yV]l
���B	{_:�gt	���X����q���	�6�t,R�������a�� �F3��I����w�i&Q�������NB�3�I-�7A?��5W�����w-��<כf|E�Ɠ�P�jU;�Ӱ�r����кg��K��s��:EWS��ƴ�6ط�Q�7�q���N^�d:r�z2/h�
}�W����J��qvqz�{x����DfL-fd�q����2�V]�؀oDy��5
����E؋�Lq&jx����޵�Z�`��Y������ �My��4�Sim��!rlr弜�x7�}����J��׍f��c\�BԮ� �ǀ����N��Vm���/��?���ܱ&`�p@`T_��w ��Uc��F�s\x��O��;��+�t�(
�;����x~'�I;agkye��A+�\���=���c�z`�)���퉡��Fr��[,c�5��YD �wӷ����5i����"��T�T�+E{mGW���C���:ݐt����}[����萪Y60h�����1�<V�/�wF�7��w��G*� F,4�S8&��
xG ��&�NP�|i�����r,Þ��hT�ص�/=�׻������۔�9}�ɏ����y��K�����rk�O�7]��W%P�V��뤜^��z��u�i��߫�/���I\�A08��t�ѫD-c1J&��I�o=���tKJ��һ��u��h�0�g)��٥�q,[����������XL�Ƚ�T�L{:�"K��C8���[Bas�����H$���|P��+���6m|��z�eI��'�*�oDDB�4~���]���-��T�S�(��Ȉ��'�߳U��3*n%rGb�^m��zND�:?G�V��H�S��֝H���p�~�p�l���O��#�)-�\�&}SEs�0�@|���
�/�#�dPSR���_К�j�Hr��%�b�-�g�~�p	�{|O��T/?m�Ǝ��A&�L\�yx�0�^��4��I:�%$��Ջ��q��Xi�-׼�pC��i��� �tt��4\�%���L���%v���	*�1��d����LR��T�^����-���O(�e���c\�z$���wW�Ǡ�/ǩ�Wiq:OC=��L{�����TH����%.��㋠���P�#Ͻ�Dpl��	�K��tg`�6I%�gN2-��$/��k���eO0���vp(����
43��Q����!����Y��D7�8�KvV�̪��;|罭�f�ߍ�l�?k�W� !��/=�C�
��^�%�h��N���_L�`�ݏ�Z�$��D���\!K�τZ�W/KS=�o�K7P�};ֿh�Xo�9M�TȬ�́d�2^�"i e/�z�p����?�J<�kZ����t�;j��xDHsi7 �ő��^%�K�.���D�5�3�L2#?��NN=5Mt�3�6�"� Umg�?S�|"���c��.��nU��|����~ʭP5�t�s�}��!�#;�d�7�_� �
��޻��/7��]\�w���c�!a�g��s���Xh��k�{����d$i�bF^����+���N��/�>X����~O��+�>���Ԏ�{�����r4VB5�I�<���=�S(��t�g�Ť�x���۲��`o�uH�~�k��G�����n1������s[#��_��0~K>L�N��g���]Ǎ ˊy�B�w��Θ��O���x�G��;a�x��Z���3�,\oM2yS�#���y��!&�sʙG��0���˿1�-������8��k~ｩ�:®��h���s�JF�H��>T؆Kc*���N�u�b9�N}����K��y'"c5�I�5�+����Ϗ��v��lZq�b�`G�Rvy79�TJ٧�P�7:���T[��d��|�7��W5~���Ӛ�h�Dk��d)��Dj��T<T�����b��e���!V��4�Ȗ&X�pp��.�2z�/�]�[tp��~�7�r��W�q�sNU�1Ƞ�k�;,�(�Y+�p�����6��]*ok��5A����!#��i`�_�/L@<�rνq[�8��b1L]	�ʘ7��#z��(y[�ab�֣G(��ϋ�ƞ{\`7D��vo��Bu`|��%g���$�CVx����5C~Z(��xF����A~8�򞳪nć+�b�{�/������X�\R���G�I��$;T�;�+K�i�-G�O<o��  ��*���t�?�{�Y��v[��9'!2+G',eX5���F�B�\�ίs�M�%�h�����r�L�c�l�i�
j�P��b%3!��z��,Yq��;�U�/�,�r�7��k;�rP���#4M�gTNb42�N^0	7yx�Ʃ��$A� I�Q�	�J-��Y�rh��by΄��>ߔZ�d�Ffڍ<pM�nP�ԇ���5J��*@�*oG`�)�V�z���f�/��7���F���'>�2���ô�Ӗ�6���2���wъ���J��?>�e��U�"x�(�3	�c��[�a�f>���Cw�NB�@*��G��wk�11�.?H�ҙ�Y~�{�h#>�Zu���xPS��O,��	���o_ɨ��d~-�DQU�|9C�����{	:(�'���K�}�'Z�K��Ѱ�C��	�a�W�F�.hEYp�P/]�^XF�|��\�����3�JloN�`��p�T:�&��ZM`"��es`G|�rHn�x(By�6�Z/8����M���#➚��'���v3�J�oA�:�����քck +���L�?��ο�1���4DTn��ߋ��*��G�Wz"����M,F'�cO� N�+��J��28��~�k�x������!�$	�-l��H�����7�8��=d¨}�>~��4G%�Y(�L`Hga�M�
�Gx���utQV*�aD����wi�?ѷ騨2xЙ�Y҂ t�8���`É4Ӻ�v�o��׾KQ�h<���l�d*�TC��L�:e�������4�Z������׎(�R#��E���lq�*D̻����j�$�q��􎃟�np���A�V��Tmm��D58 �S�;mL��՟b!�{_1�(�D!�m��~Lgem� �B�#�2��R��e�f4��{�g{���&�\.���TK��	EM��^L�Z�o���W�-ѕT<�_��L���W�=4�ӂX>��� ��!烣��AE5�+-�n)�]'�OO¤�����hTٗ��
R8�z���>l��Մf��Ly7��j�B��r�Y:��j�L.�����׳��+��<>5����i�X��ܸ=�m,'����<?�*.d 8,��j(�#�B�5����	^ih[e��-��ې�ca��H������;�PfU�F,)xӘ��ϳ�9RU�}i]�jS�����ŀ�
��q�
c"˰��ar��h:Sq8�)o�����~"��a�أ:��:�:�_J"�]��K[��	�^��Y�S���߻��x�މ,��]%0�%d����T�����)�w��|��������ო<�,(���e樿1�p<+ڌ��H^�DYY��E��L�߈��h�!�G1a��� ir���3��"�����jGr�[_��y��hVSX����v�NF3 �-p�)#H��8"�����j�qV/�ʄV�|���&8� �J耴/6�a4�'"C��ƣ�0�f1忳�G�E�y[�7Rq�Ot����̜+�/��rUT���C�����1��܏�Ƒ�����=-�xz��e�x�-�qԶ$'B٘��!�q���JAY�5�;��IB��%��G{_�2��Ho'KK21�B���׭F����ꌋ�e�P�&ɭ�"����`C�W=k��8w�V5�7�ȶw,���\�n8��a`�2���!�R��m�c�+�<Lp��?�6]���M�Mç�l�2�I����|L<|F:?Z2���}�����3����"B�	!�.D0�M�`�q���:�"��ZX��K�W~r���wg՜���La;g�:����Z���l����E]��T@�v�m�x1�E�O�V�/�HZ9�]��5`��If�OqE:)���E�dl�����(
a��v1/@� ����;��acw`�9*(w�p����Nn�䮁�#�>*��3O�L�����旲�T� �g��{�� Rژ�	~w���vO]�> Q刏� �W��j��?��"yȬ�$�V�\��l
�٬���M 0�b=xE0�����)m�;�_�ݦ�� ����-�#��B�*O˿���,O��_��v�Α"J�p9 d)���w�n<@�{�����t�ܤ��S����c��d��=�u@��BPb�����F_���p(;�$�d`���L>�Z±M��d$��q�r�=	�:7o�"��ˬ)�z��2�&��d��$�=Ķ8k0�(�B�D�����h��C������Ow=�J}�4J���w�p�7�ĘtV�bY�`�3Ƙ��G!� .���&�@��S�0֛�p+����6��O�c��6D+7w5c;�
�o)���%oI��'�*צ�q�(�PS �Э���>7�O3<�9�Cq(z��-l8���?F�r�	w[G_�h+�/��7(�&otx�I��D:�}��r���D�*��ڔ2�$������n�Ɔ�\���&u�0HZyzE]�C�U�o�hq�YH�1�_'9�Ӿu��_G��`~�tjS�Sa���3���3rF�ʇ������8���2,j��>lfv�)�Y	Q�*k����r?�B�.k��:�%���~��`�C�B�ܱ�@hD:������dd�O�F
Iw�z��	B(��7�J�����$�ӻ�t����rtF3׍�?�7[\���2aƶ�Ș�>�5?k��j���pnc�1e�k8 t�=�Ov絏��w��f�Wi��f�̙�,�)�!;k���q�Uɬ��D
�*
9Ύ>�-�O����	��Ǖ+K���2���'y>p5��j�����[gk4��ϓ����3�Gn�G"���Q�Nٝ������x��.~�:���0׸4b;	X��{��0����9'�N!RxDƅ}��IΏ���y�,{�
;���U���EjE�MH��{�t�>*�lr!e3%H�^3�8�ޚç�:_����-kX�|��ef; �n}�z:6�bj��%��r��1,iyEA�b�}��M1~KT����W��L�B^�����+0��<�UC�:'"%t0���Xo�"h��0����V�/��ju��^4����<Es�t��]�u�".&��x|�XA|E;��v$~4�~ 	����)ZO���
�=5N�X�ݩױ0�Q`����Gɠ&��R�F�-/v4���_4��#�:��ay#,����M" Fh�Ґ;fb&�Dƻp�
��?�� (�	�&�?HkN8�������(M�L3J(j|���pUO�����)�-��_tE��S�Mb��E�P
� ����!��$0r(�2������?OJN���AT��Q��"a�-���I]f���Vu�ď������nڤI�=��;�tW����SB�*��U�
w�IMl���u�'��L��>2�\��A��������[�W���#�s�ڤB�-U��!.���!����#�;%���O�kL��]O]g�pZ���ɹ�M.�U�Y�����s"e�zAvAL��R���y�ZB�$q?�+~���pޓ�eN�&8T�`��'�L�Ȟ����UT2g]��'�6�r���#w%��EL}oUtf��L�=�#��+ڟ���p|/���>���M3}�B�">�=��[kE�=������&���~�==31�Z��m�k8F��l�(T���_���n��|t]��s��I�E�)F�\h��g�59������[}�Y^��D� ݆|�"�ͽ��z֩����F������jY
��[00�so!��a����AQA����j6c�RT�����\���>���.Ix2
\�L?Y��p1�
������9��B�^��+��� 
���J��<�������E,�MV%'>kZd�z��j�����c�l��x���y�>��|���ΎFCI��c��S��"ae����Z.9� �*�_T]����wn��98�)����MƂ+��
���Qk!r	f��uu݄�y����v�fՀ�ʃ��X�0��������+ɕ��Es��;��Z6��M�3'��a�N#�X��쀑�<�D��9-��C�Y%�u�h�ʜ:�D��i��	�!����T�x�5~s2w�C��voIQ��.�����&ج[������b�.�qʛW���s���G����K��3�ܥS���E�v-�~�9>���=S+�U�7֮+>�Գp*�h;�$���3~�(;���w���Ճ��c��H�Ib�]1�[��F$�G�lwp�͉*���Sѹ�fm�ǆ�������i�+��Ks��,(�n@V>ۤ@�̃�fK�ɴ��޵0���@�� x�-�-b���\��~�-�����b^��C��V��u��{�_:�srz!C�[Y�}��Y��r���"�A�y'+���8?�{���ٳ�Gr'Qg6�q]��w} �B��OSe�1Sr�&�=�î����{PA
�
�:�M8_��'�������F�o�<E0��<LSR�Y��כO���F�or�s��0p����XH�y�'nTSP����[_�K[`�����/���3@s���C���h89��+(�@�o�Ez��W��ǜ�p�M�\�qvz#��Z��Y��7N|%v�+e�G����Y����C����_�^�=uCKK���l^k�Ӹ�,��7���~�b�v/�m�l�����a��{1�ܾ#Q��',B������KDH��_�p��wEs��?��|����렣�h����٢�u��&	�

����oCԲW%���"�������"nq��;TҪ�o�Bڀ�9)�}�T��u�*|��]|>(�� |��$R��G���㰷o���V�`�-{L'
k�nz�������U4p������R�����kPYM�R��b�G�8s�lM2	���]�����I��#�Z���qR�ﴄZ���n�L34wn"��B[��W�A{mWx�.�_~��>"a�iQ�*�!4�`��U%�8�	��y�v��=F�����h����bCKP��/X�(��(��:"!���	�M�i�OY}A�,S��hȿvRQ����J���zXO�X�8�^��t�J�ӭ�L�d�ݵ��F�2G�g[����R�O˫H��ƫ�3ny쬒�g$�Y��XS���rgƥ�i@���
����+�-�S�Q��"��V1h��C��Dr��hZ69M�t�S
4e#��$�ĳ����sM��D���k�7[�d�'0���젥Cm��
�K� �E�R������0
���p�N���rB�-5�⇳� tc(v��ݹDX�} m?���8����I���"�a�����7�o�l���9�	�O�ƗS݂��M��%�����N�E�Fz$�õ��*z�t����8T!�}�z��,n��Zv��~�]����92k���z}��c���~~��`�V Ԥ��Ѣ�4���I��F��g��aل�qg?ѵ����b�^)�,خ�����|݈�U��JK�����u�c�#U�5E���/�q�+E��1ە��8����4
�����0Z� �.�"L�*����c�K�I`{�<QE�r-~fٖ�'���տ�r+�n���=�I ����7P���?��y.(\���a��b�n9����^�7B���sm�@_H�MƔ#*��
�f��^�l�sS��Op��׭� �	��8>��=�ȓQ_ؒ���9�n�K��aU��]<e@ےn=ר)�9����s�=d�!���?{��||o����@�-����郂6V��ew{��Ϊ�+�p�񵍎3���X�a?�C���WWW��L��AA����[�q�X����Gvb����C�A��?jnA��6��L���<����/���j�W�^_���߳Gf��D�U�,}�#�g`dۮ)z|E�<Ti��u(Q����`�� �,9��IiԼ^t?�\ٳ�2��̕4����N���͉��{��=G|H���l�Vۡ0v~oI�
p��y��U����F�VFI1�^���ŧ|����6�'���ޓ�b�98���qM�T�%�e����g�&��g���/c^L����W��]Y_�������hg�
� a.&��%d�qvF�UK�m��G��(�ix�����x Î�	�+I]��r\���@ŧ+�Du{����T�p�{� �p͟)�q�I�& |�T���34�I� �C!C�!�=�y)P�D3��C?0x�,��W�7#B�|6D4����7PB 3�Xt#���Z�� V�N�� �~ �I}��l5��-?q�O���~zz`U��!��*a��̍M?��(u���f�M�c��#1w2���_�x�\:��(�jfs@c����M	x~�RM#�Ҕl2]F<�^��z�0}��ٌy�Ώs���(�@�6z��3/I����mY�����l@2����W��6n�%��y2���s�O�ki��-���M�$K/�aI�&(�Y�bg��ĉI�u����,r�s�}�X�5�v.�?qF�w�J�33�SC�\n���la�ZM"L��֤��O�,FxT�I)D3j���&��n�ZEEuh���6��W&�v��G����f����G���l�g1�
xE���(V	
����Mm}n�9�l8 �=�{GFa	�ѵ�wd`����p��?Z]��_#��OG�E��	�u���Җ2�;��nN����k�ȡl���<�
�*畐6���|}Yr�t��]�|�,���^k��E�KE�xdʗ���P���Nv%\�F�8����h�����@L�����F���؄^И?��&1�>@�r�u������T��\�9��!�7I%w�'Bx�M��^�]*�7?�'m��˿�6����@j�*���v��)(Q�	<(m��m��W�j91i]}�,�UI�_ǉ�=�?��.�y�7L-V}�*fT�Uvl��^{��N�ڸ{#ꂫ)��)e��f����p�{T
a�a�k~���j�;$D�:~�l���(�֌?_�6���0���_Kn������1��]M4ދ���0u��7��g*D�(H��F��h�C�P�X\f|�j��_,�5����O��t���[�> ���;98y��j����q��+���l�;�[������ލ���	��L�`҅����]�����15�$K?E9�D�ÚS�l�hl�i$���볍�0&��,d�3 V��^Xk�D�m{�e!+D/<=�}��b}M�c	��lr线jU���]._�D��?�x�G8��α�7��Df����8�%F���3RA�q�ųܩ@��L�z� �1��!��s�����K�󣤨$M��qEߋ<2W0Q�ơz_�>�Z=�;����jA�MSRM����݂!��Oi���H��0�BA\lw�4z�{9Ռ�6He�O��{��n��u�=�UI�s��TB����+U��y%��N+`�zvQ!#�PH �!�O[��J���?&Q���8�l>|7_p�����a �7ha�g��;۴�de5���,B�d�g���
g��6,�F�gNJxD�`w�%�A���	�g��g� ��Q��`uO΂*hņ9^��A�l�MdҀ�[%p]Oש!G�6�Y?H����$��S�P�u�p�x�#OLE链#{[

��X���i�_���U�'>�H�2L�����U���a��<����ѻ�����>�6��k	-!�n�L��� �f�t(�@O��pD���lB�or;�Taa�GY^���59(�a�VI�w����2��ߍJԕ��4��	�z�rWh����N}<�W�����#<6�XG��}1���;$�z_F�K"�e�ˊ"������~6�+��l.��l"q��bl�Y�"Ӭ�o��@L)�mFD� �����(@�幠(�O[�Н RIȱ��_�:����;ȎO��l�4Q�"��`3ԇ%�
ne�E�'�A.���(�嫤���.�Y��B"�XQl ��'8�@FB��I9 ���
<��$�x�<]B��<���Zďp�����������ז�U��T��Y�m�):�
����;!A��,����=�(/\��2��)���o\����o$?�<N�9�8��ab�Dz��	M
JM`I�3,q��C�"k�~�zB���:�brz�:c��UN��kr9��fJ��Gd9���biZi%������p�6�����[��j?M��n�u\��3Bhit4h��=�N�8f��N�����ឪC&KP�05Ӭ2`\��ħ��;�<�3T�h1���w�@YՃ"9��x����o�wE�89��M�k�t.M�p ж��'(�֨�ok�x�~�f��4�uϺ}6՛aͦ��WX��ࡏz��)}�D.y�$Z	m<ԟ�'��*,䣟�����f�Y�J&���3��P�в�J%g���3��&�!}��i��f[a{�y��ox��>ۇ��+�F�� �M�͑�M,SS:ː�g�۵��!�e�d���� ���N8�c^���@�P�o�g���@�}�g�"R���?kN��?�1ﾖ� �:����] d�����J�3���#�����
�8�#0����/���q�����=}�]��+$��4�Xy<���73���B�)QZ�OtS����xc�s���m�HJ�l+�T���B�4���CT47vO"�<������ s�AG�xR^t��e�v	7�;ƒ�E	����m� �����vEٞq~�̽����T��B��Y���W���!�)���!e�7�
���p:�Z�Q�Ǯ�.Ī;*��g?��%~����f�¼��xac��|�h���|�Ϳ�Ա�)S�eo��JdPP.�}�K���|qǊ��U} F�z#Á9���Q�O��""b����d��!��g��6c�I!�^�	D�H2�7yv#�|���V;6�w R]C�U}J ��p��w�,����:l2�2��M�0!yݬ-�ϥ�;�i��Z�$�&��[��8�K�2 ��a.�At �^?�>��&���I:8�:L�!�{�Ҕ&��A�̷�2�&�E�Y��fN�>h8�Y3�4�(<:���"_���-����A��y����<'U�x��+��bW�&�� �
�wz;�º_N�0������ ��^ w.��L��k�у#Z�5*�KWXy��<��x��x���������%~����G~�q�M,T�T�-o�C�'�E A�&�Ǐg^�kP�=Q�)}�Ҥ�f���eMs%b[�]<S��{I+���ۂ���(>����փ�����Bw�����į���x6�k��}����H�,��P���υ�"g܋���I�Y'��w�.�f�2���f�2�ep�p3�ʐvE��3���ԕa�~;�B�Xpy|�̬�JgO�8��l82�ތ*��)c5��h��tbQӁ�pf�^C�[^s�Ь�����D=�`��<�;�������y��CϊI���,d���\@��1�!�ݱ�!���X�ޠ�	�@E�-��W��.�|ٔ�'ՠ|�h=<��s�_��(�i��w����7�|03�Rx���͓Rb�1�!�����U?r�{�hO�N'��t1�*�2=��C�9���U��84�ig|	̍��\�
E�%�n��ZuB�j����b�pN��U���?Rh�@J1<�Y�O?��XR�⺣�G,,�Dr��';���;��O��7�	}�z[�����U.��5�̳5��P��M�����<��[��`&1�S�5SO`�T�Ё5�ޛ��@�'��������g`��Ϟ�sQ #�������u%���f~���]z.<����0�1q=_�a���T�����A����yy_g:0zCsX�o�P��iҮ����ݜL�uM�}���A@���mʻ�ޞ��j�q��.�-�w?�ݎ����b�v��RЉ���hv&�Q{uC�C�F�݇nҝE\�J������f�kR��-ش�"�
�����W2w��$`v]�1!/I�(�5�s)fB�%~��?�ER1h����X�~�[���>v:�^��%[�ʀ"g.���6 �K�a�HXnP�sS�����}ϒ!H^���?�Nɔ���� �*�KIɰ� :��Ԉl���O6�ՠeQ:�e�?�p1�Zm⮏����<b�/݁��<H��e�y
N���)���z��`0Z�/�.�v����׵�m6�exB<�k��byn�ɟ�v�=e���������̹��z��z2)�^����3Wh�D�
:��'k�6#�N��2 d�����5�!Yx��.���� ��zSA������Ll���M�4�@���|x&������z�v�Rr��ַ�5h펵F��eAqp�|&��\+q�	H{�Q�jۑ�h�x�o wZ9`����_5�L�sIn/ѿ<:8� R��к�+\�F���|0ei� �P���n��QXY�x&��5.H	=����^�B�E8�HNtQ����XK?/#ǭ����x�,��ى`�b#I�2�(o���=�W]H�MI:S�=	�\���M{�]�e;�?�-�Q0�<6`
_.���3�A 'I ���&�/��Kc2�E�e
���3��z�kc]	 ��oz����q�f;�K�T�Z(-r�e�p��oH./{D�<P��6r�գ_���&����Zט�J��������ě��5�䙃�H�ZY���<��ۺH�;T�<= ���7aɆvͤ��k�����Y�~����K���.�q3���[�hˬIZ�.xb�.Z��^�K��z���g#�rxD����6�P����L��h�qe���>d�����n�T&7B���ƃm�		hI����@a�K1�@ᢇ	�+��`՝���Je]����4K�Ͻ���P��-��/�<���d���*�]5��w(��L��-/�ZҦ��^�Җ �����{��̓��Zz��3$7�8{�5 �K4�\��k@M�D����>��!nܺnD�C�/�3����]!|B��8><��R�gLL�����*׺�h���O ��=���sǩGC�̷_�E54�vNK9s�ze�K"jF�@3�5l@��h�`��.���$+��)v���h>�y��z���f�S
>���#�I�Z���Zw!��[3�`�Y8��<�<Pbw��]��hk�建>�i�"Y���cG�b+��9��a�]`��i����3
@yA#���2�����Q$A[����#�o<�֛��I	�E}���_ۨSZ�vDI[H$2���\�<7W"B��`��1���"���(�t��*���[��dE��-�vS��
���?10�LR�٫b��Tq�'���}����]�Z;jL�.��zI*C���`+cg��� �Ht\F�ie�.�v�,ou��`B�&-�rd�	!�,�f�j��������k�j[&!��l�� a���%w{,..�.x�lگ�^_dy|W}������l��d�*�'�:cu3�{��E�!X��LJ��9�0� $?���0����%���q�1M ��X��[A�߿�*n�ev�3Gqݚt��ނ��q^3�a}�M|Q�Y��P0ɘg�I�4KjIQȊ��2xoo���һ6��I�}`r�,��9.}B��pܵ���
���JPa�Z��q׃%���kш���8����|xf%�T�i%�T�;GI$i��ެ�LgĮtt��Tޞ{��A���u1t�!��@�y2;�M�"e�jZ����d�X��z/5x?��!\�ox�v��.��!� �G�[zk[51��i�5gF���U�d�y[Z����)�~$����G�v��֕wD'3���ˊ��i ��G�ͨ���r#%-���Ǖ�l^��L�Y���"l�%�+\���Pᵊ"�ԙޮ�*qI�h�08���h}�1e�7^<i�p=�@�X������BJ%�h8�~�<�w�>	J�[^��>U6'³�甋%ꠋ���m��~��KΙ��o��;m7�P�o��:<"�~�_�mTk����C/��v����h��f�Q7����®c���T��n�<�j��7z��*�`ChJ��fy�uC����Z�wH=8�H��Sw�j0�!P5{ۄi%Ĕ�̎ų$��\��-r�/�b*X3]��ׁ��3d��5� �Q�Y	�5T��F_C���r�N_G{����=3�\�}��6��e�f=#��aBqM���9�$ܨ��2�����L�p�*���$rm<�Yj#���T��W;u��2pwa��(#�| �1����d�R���0΢����V�NQF���өz��nϹz˒6�zT6,��18Zؘ�z���wT�t��&���Zx�A��}S0@e$�$�Ӭ�O :ȓ*��I^��o��<ͫ���F{_�!*��*��"AW�4�j(��L����'%��ڪ��d��0ڻ��=!�FWlv9���@m�.�P�ƀK�W�1�ۥ�� �=(Z-�J�I�����'V�	&~X������W)4;W�O_Ⱥ���4G輦Ic�b̞�>�J!v�S���2<D�+I{Rfd2�)�ϛt�}ܑ�Ѝ�zi�4mU�pd�F[�:��b���\p$�WX5Q�<�g(�0v85�?&~�S�g�t�����R,���!4/��:�]�� O�`��Xk^&���*��."�~�,�	r�|.M���1��՛6TM�~M7��5� cf�)�.�E���G1��.�+yւl�ܟ� ��������vQ��b����1�������j�V�4��%�h�<�-j����:Z�9�A�
��:��,�
�,^�rϴaV�C(7&"��vl�%$Dl���e����_\o�o���*:k��+��U:x�꺻�*}�B_��q�P�[B� _�&����?གྷ�\���N9��n����:�u��%��v)�H�.ML�R���%MT����c���&��;`��@����}������R+m�s��Bo`��<�l"�v)���{!!ַ'I}�YEsq�ElϘ�a�]M�ǷN�;�q�R?]������l�/�	��I��>%r_��b���t�g��1���4�bΊ`��8��x����8���U��@�}}�;��g��꬧,7��A`YJ�;�ͻeJߌ+���$\#II顭f����z�c��o �L���(
�8w�xE��R��4O{����/K�l"�C��P.�ȋ>��8������J��i�7%c/>~?"�I�C��x��l������Wș�R�cOظ�_�C<�6Y���F�?�=�Xg\�e�!�*�JQg���#�u�������Gȋ|h0g����ם+ڸ��Ӭb�Í���r��:�\�ֲ02�4��]�$�ծ3-c>��K�Ы�c.-�9��}#�����|���%�_���s9����u[	yfm�	^ܾ�H����%{ṃr�����&��!w��������
8�'����}��k<��t��#`�;Yo�9뛄i	��dS���ML�YSRag�Đ~*�(&�~$�eh0�W4V �6�������G��s:�{����L{�OA)� ���ʎ�^���Η5��Wl�Qs[!@	AF��Hz���،�?��Eִ�,F▼� �|OL`A�U<�%չ�K���j�IQpN�:�-S-�|u^I���8M� @�����[�C��{���l� �"�]q�6������2Q2��
~�,��F��e�N��eZmD���M�j���_�����O���Q�b]�8G�HW�~���F�N�7��^�[z�4I��Vn�&6%�O��~��kW��p���#������ߨ=�;�M���O��
�F�\�-z�r���kAl_���9U!��:�I�I����is  ~&%)#/����gd�P�֋:A����?�D���+�|�*U��././Yq��p�@F���s�a2o�<��4��jѯ���EkT
�����jGNo*6JS9��c��^/ɂ}�(�,ȯ����)k�������m�7�k�. �o�έ���-&�:I��2^�-�K��q2hG��Tj�M���b����j����,�J|{-<��-}r>D%Ɵ��kuuHL;>=0ґ �d��Ώ���%V��0��Pnov4Ͷ�������>��%~<u9?V9X��6�q�� x3�Q#����ڐ!��ɽ���[U�V�x��`$�;\�ٞR��k���'��y>�ɕ �3���ڏ+�/e��'���f���t\��Ջ�����'bEuД �$T7��`��uӼ/ ��IУ�������}�Ŝl�Z��?ڮq$�  �L�1$幃����lWH:|CA��ͅ�z�]�d�3�k�N��a��?#����� ��~p�)oD���ol]�P�(HP6ı�P-�����q�y����r�V��%n���b�����
ǡX�V�.=���zk���2UhqD�p��j=�=���6u�vY�P��!�d�@�G�9("�CY���h��@�z�wD���)߅�X)�F1��0�ϹYh0��|8 ��Y�L텯�������SS��.b���uR���G�7W� �BBV`ĭ#7��-4t�A���ZWB~�.��W���X �+-��W��*_�Ir��FK��{�]�8VG��o��$60۠���ϫ~�aWYDtj�,�$�ɪ�ܧ��zz�Hc2V^�0<�J����i'�Qt2Q�jM�H����C�|�ڬj٭!Of\.�g%љ	?&CFمI#�q���wg��$Ӑeg�����`QApۍF����kE��(���^��o�����ܲa*�9��sf>]_�����"���T$
�<)�S��h� w��Ӡ$ȁ���t�ޣ뉫��y��x���}�����z�>��ʮ"����'��q�@o2�-�8�"��D���*����Ѡ�r�d�{V���Z��b��5����;3��.��~䏰�;���-�� �	Z��'�:N�
��ȫ�+�jZ�RY�+59�)��t�/=~p.x���� �rm�B[�6��ձ��s�JH��+�
�v��$���P�-�9�:;�Q�E)$�t��.�z����N��Y��쎒� ��+yX�?��T���?�Ӱ���$�y�F�;�A����1����>Bv�=$!;��7�u��5�Ia[�+iur��X4��Pފ����o�*�,���T���#�eB��<��,Ӓ�}9
�#PJ��P�=]����uʻ��z�U��K&G��z<���V���j8����� Vy��Mi�̻�:4�"�b$n,�0�y�%�?�2:?��Ji�^"q8�[�![:���9WD�k	v��ߩ�;�A��(QI�"�dɀ��K#��u�\���L>ʧX�^"��`?��7�\\ �j%M�����O	�IL�l�dZgJ���1��Ւ=h�-��bX���fݻ!iԀ�y%���D_4�޷͒�`Z~�mqD�x�}��R���R��,J	!7	�;��!us+ 1J^�K�v�3�<3�T�<���il�O��-N	���J��������:P�p�����hS!�O9ً��3W�i��1�R^��4�����1�Xjv���{`�egx�M8�h�w�;}�D�5C�M��(b��]~cT#X�wט	�l�׏y��Ѽ���X��)�G`0d���y�|���#Vgӗ��{��������t?������g6.���:�%��*$��gIv/g1��iQ���p8����x$B�9����Hu,4��|��98��Aeql`�6��MK��Ii)�yY����nS�G�������F�j�hBf� P��:�"�Q4A0[�ù���;V [(��@V�S8�&��G!}Ί÷t*
9�ͣ��;��ֽ��쎊Þ2~:8��B�4�r-���L�@hH���J1��2K�0va\�p�_��U-1/;�hHh;x���w�w{O/z}�Z�ڡ=)u����;�A��q%�/�����2Nj�\��b�i��R���K�^"�b�`�Zng;�j�)q���T�s�S�ud�C��y���
k��4� ���zF4��~��:$`�F�nS�L����OetE#����J�w�y!���W �����ѥ�.=
�_N�Ip76�14��M [d;:��q�o���g
@ϦŔJ?�KK\"�' �V�?t$����M���i�j��@٧ot����9�ָ��gئw����cI�2�� 9���X~���T˸N�q�A�����zW��� sqt�� JA�t��Q%����n��5~������(P�|�G��#b�� �ky��k�_�2�c�C��[Y�f����J3E���<%1g:�'>��������0w�� %0�ռ(�Ǻ���b�[�ђCr���@J�?kD��,'���F(�m��Rz�*�ґ8%ǧvR��X�����y�YO��a�WX� �(���`��<����ď�9�r:�y1	��=���0/Kch�-L��<�_7D	�a*�d���X���1#��b�U��}�L�� �#G^�%�4���H���bZ���Ge�µ?o��Эbƣ��_���g�&����v�gov�Ԥ�ۢ0�6V�\��g"j�PWb�ؓVYXT��mb�������
�.j/�<j3Z�tF��uy\*�Aa�I;9�}e���_�;΄���X^H'���^M4������6�!'� �)ۘ���H���nTwRt_��4h#�5"4GN=�A<؟\�y5�B/e�}��Mx��{���j�q��Q8�v ��+q��9����0�U��$g�Z�"ָi�j�>�Bu�ڑ�::=�`eR��]�r5F�-t����[�������!��9�*��2z*�����>O�9�=���E��Ȏ�[�'?�9D�|��8��D}����?'Q�,:j��O����5���9p,[�;M橌J�r�v������d��6���Ĥ�I�}�
�'q�t󗴀�\^��E��P��zS�,p&��Ӧ��0e���7mZ��q}5��؎u��Ex�gJ�m� )�p�@�g/�	_}L#��f��F���5!�4�-O���"��F����I�����v(�׮��:�秢/?�礽����s��5���I1<���3+v ��8-0!\��#��@{�CH�&�����Z=���XƤ���o)�3`�Ѹ��"����ϥ�,A���
���׹2�T=Fָ�����8����I'v����O�|,��߸Z������OUX���'����Fp[�l'����-�gw�S��N�y:����i�稂�����S|x��������`;dᡧTX�k/��e���Ns��<,��"?&�}��G�W�����i���rZ�����D�~��v�e��`�F�i�_hp�v��;�~Kl����>��h��Z�q1p^�a���Ǝ.�����m�'�:��В�y�6$9Nf�3݄T-����� �W_xÑ9�Ғ>׉6z�c�|,�	F�>S�1-h7��g�9Y4�g���0�	2<�3���G��-w���-������Z����3��8�X$bH����M���9��b�@|����Xxn�91�����ܪ�`�]�k�YC<��63쟹6ӮE������e*�C�?'��.7M�l��?�O���q%��A�^^�����l�E�Y�ԕd<�ԥ�[�8]���"���0"��)ػ���t��L��4��k%>$$Q}���PG����{NA_X��_��o�`���vL8 =� *e�����;5��:<�L0X,m3}��	;�x(����ݣf5Я�=����|��9�*U�+�n�e~��Դ6Q�A�L�X�:�I�x��4.�[�2�p. � ?)��Q���g��<N�JԐ�(u����0�uk"'���˕�Ra-�Z��R:��9�D�kc0_�LMn��)�tPֽ	��9�;�m�^�$������B9.ŗ͗hm�ƿ� h�F�q��*Q.�b��`baL>��Seyޜ����"�]�ddr����:�R�����Z~����Z�Ni��yB4&*��i��=�f#�@��WOnu���E����r�}z�T�|"])�b��U(�)E��5N��O"��:0^0�V
xٮA�C/��2��u.�'h�7�ӣx�׸_a�^;*��˓�(�P9o3��VD���	�rK$�������r����af�豣PS�zi���i/P��$@���2B���q߰ux{I��8�"=�fZ���!k�ݷ3�F�G��+g	���U�0�@Uf��}Xbez�����,@�w�dw궤q��`����7�����yp'V��cR��ht�uwע���}�y<�v���呛 F�H���_��5��|x�ӗ�2����μ�"2<?�l*��0�.�)E�g2�h51�na&��-�=��fG�Ic19��{� '����<l�839�P��\2�=$�d�|	��s����*-Iw]t�!��Bw�W��ء`an��qk���o�e�V;|�Kv_,�Q;@�;��������=�o_e��j�`�N��>WƯ���~�kX�r#�l���=���s��`����	"��/�$7:�e{���G��t�^X>:95������i����W�`,�W���8����m�Ro��`ۥ�:x���2��ОI�x�k�>����v�<���_��r�����Qݵ֩�(���I �@�4��=��^��YH�Cj�=�h�����E$��!��a�DQjT ���y�u�@���M��0�=|+�c�>ִލ�H�������g�)y8�ׅ~�d1�oEu��k$�)O�O��K&���H?����v�W�P�:�|-���8	����;�-�V��i��-c�h��R���KSH����ŧ셏!�P
�Ƒ����o���<�/��<;̚iU�����[ѭh^X�b�]�<P��+���*U�ҁR�V����ݿ<����d>߽r��X,�7��?M��!��@�e�EC��G�w�57��^���)Ls;I�<�y-�YI�-�f��g�=j��=�eaO$z�q��U��F�޵�pQ�<pm��f�<�q�s���X�NL��K"��>��o8Л~���B���������J���}� ��22M _���.�j���y�����m���a��M8"\"{��K�($����N�눘\>gc�"؈�(^���XRf�o�""��L�V�w�UE�ﻆ\�$V��-��˘L�\�$���P1��4�"��=1�]v�geA�]�e���+`=���0��-�}�;�[bT{Z�s�K������c�4O��t����"ؼ����I��fv�)j���ʓ��>��;��p{��J�� ��X"�Q6NP@0VIO��rk4��������<�DN7aB�q��;.2B�3J���2�����D�����ۖ�9���j��x1ٰ?G�)|ie���_k߁�{^��R�ںS���b�) ���m�fo�ϒ�-;��&3;&?3uw����
�ߘ��x����A����-��~�6�IH/VDܪ��~O�a[�k��'��Qa[����	�G�-��A����/�79�jݗ�0�UT)E��-F�H�0N\{/��D��GR���6Sz����*��(����x��a!�n�O�ʱ�b�)��P!�8�c�{]d�2�̠{�A�?���]�^\H���am[�}��\��&a��!�6��.wPsa�ߍ\v��7�\�;@+_�߉e��Cњ�n�6y�M���i��/��xW��JK���$w�-kX*?��Ę;jI *�t��?+��E� p/��v�x~;��1AϏ�:��$?7��jh)��&Aw��I�������m��Q�x����A�S�kno�2iu"����Z��J"w��m��21��/�A�{�uz�����5FLQ�yMS���t�"6hG���k1M_Ĺ@����?	q5f��!�	% R�u��1a������o�w�3(4\Լ�9A��cj}�8�ɪ���=�}��M�
����-qP��)�H�e��b���4�-tK���#��ߔF��=�-vX�W�^9>���^rӐ��4���VOw�� Tb@�G�4�py#�(>�O{��S~!G�}7��ˎ��� ��U~x�r]��&�U��H�&S���0�Iǖ���e��6VI��W�! �~S����}���#}{��?!U�����q%��s�}r�TzR}U�'��Ǚ�Y�_ҷ�s:�����t�H��
�?�Fbn0v�3I@��a|Ȝ��֣8�mm��ZW�i�x���.M֡�q�NZ;W�*�=�-�S�����,�V�q�U�A�s�dg�YD⡫2Hy!C�M���/��S����%N��Y���x�CF��k�>��0�?�KPr�TX��gj��!,�f?��:wq�U~�M\Y�AZ3$��x�:9?�/���t�}E�Q�A�m#m����	�HO,�0yDz���:I��e,��zh]q����ں�7�t�%`s�@5�}��~����{�kx?��te�I��X�+u���;�z�-��=��n��������R�D3����Ș��(��L�JF�k4 W�ס,�k���{o�i�'S�xؙsy�,:X[��)lv�����yT!�v�ưɕ��̺T��눬-�T�3t�1I�Ad?�@]��9�!	&�=y+�4�:�ccO(����[�s��Zό�	\���}q�?�%�9��if��Sx�@��F�}u,�.d�Y��l��ƾ�#�ˋ6��;:K��*kJ���Q��t+����4��y^g�|1̜���1s���_���~a&9�vD�ճ�������sLM����÷JED�ץ7N�CT�<���%\�d29vq6ΝD�`뀚T1�Δ/^Ei7�+`��>eˢ�T���v+���U�{�8�{\+j�LX�LZ�#p5��~�(�D�r!�]"��;Z٨~p��!s�"'[u�Ww���)lXBz������i����g=�����7Vs�㜽1���T�;]�/
���#���C9עۣ&_���N�o(`û�zo�*�_5�t��oDG�+Sޘv���
I�����JX�M<�~(���!��+�@�՝�����Z�D���h���^	a����L��X
�X����^��	��%�>X�i9C�]\#j�Ș@�n�x��@*�,8@73���´�&�6��4�:?#������Ϫz�I��٥��;�ϤH�������){����,���MoH�S<�����X[��$�Ƌo����.�8���A-�e��g��������%�&ʈC��ָ� ������뮘|���J�d4;�׭Y�/h���N��Y�jijB�9�� ��R��
���jN�P�km�������?�j#�����j0��0Uxș41ӕ`mr*��w�!�����q(�_�7O�m�2���I��̱N1/6R8g$з��K����7�Y/EOу�|8�@��C�\�k�'cZ��r��L�0Fo_`et���J@®��'0qt�wAqU�I^�;.�gP���Hi{��Ŗl�)V돤4+�/O��|�L�`�G&b62�|5 ��،$���z�|b�{ţ ��U��x;�a��/��0Z�u��1?��į.	��Û��u~��T>赐����Oj�T������>G��Lo�8F���Z./�G��RV�����j�M��#�������6<kX�򂴫��.m�%s��u0�A�����8PJ �Mr�4K��	���m��;qs5Xp��>g��t&��y���2lL}�D��J�١d (�_�Y��P��6u�:�� ��4F=��7m^��´�I��K�Z��d��\s��:��"����:��ٙ���Lq
�zDX,�{��5��N�
��ʐ�G�Q�7X	~��.[�7�mr����@]v��ps��P3y��G�< �E �ZՖ��a�ŗb����6��̾��2��:�"8��䠻;�c7�Z���pv�z9ѐW��u,�پ��I����UW%��˼�Yg�/׹�"�h�cis�n
:n�!Xx�̩��˄N;Ϊ^<�ڳd�0[E�U����SX��-͈��usz��nZq�����Y�(�<�I�e��ܳ����b��f�W����v���N��G�`,Y#~՗d�8��5`tw�c�c݁�7����ӾL���V��/�?^Os��!�p�_#�3QE'P��Ҫ��t�]����t���E-�bJfrH����‹Ak�՝�7�R��t�.����oB������Kil�ap�h�a���n�	���rh���Z!8Ņqh�fUF3���cd��آ�E���U���1��[���+!��Or��!l�I4��K	h���hɳ�NH2���6�>�%��l��sx9^�D[��LI�	�}���fjڥ0` ��)Z6����l8!�&��nX�[㋦[ T��%|��'�b+�S�9aR�緐���_�e�N\�|H�7X���GC
Cۂr9�ÉVD�fU#	X0U�/����pU?X`S�!�-t�@
<�<�с�/�yC����|<X�����ܡ�-�@�ߝMƚ�\��c(��(ߋ�,uQ�l7Mf��^P�&�c�~���?_����H��όw{9�~6�j��˕�=��TC�o��,��鿔;��Y�(r��Xp��|�
*2YX���
�S��E!�H�@r9(�6,���JQ�@���+�σ�H�5Z2��,�*7�j�i�Zy���L��T��� wRM����|d�Ӧ�X��Q�{��b��L|f���֜�%MI���r �#k�a*:ǡ?}�I�=��Q�^X������ݹ�մ���W�N���	���*m<+�.Q�W�>�9�9����g 0�6�\m0�!���2��4�s*�[m�D�p/���#����}�Ww�
�8���V�\��������:��,�� T<�z�9����@g�8�>��oX���Äu�dF����b� �\��p�#��f�]8�眩{J��N��sh��[�|�4#��s�xt�x�J,ѭ��Ch�Ŕ�>���CP��(�K-������؂�wT+)6x�ڰ����kԗ�@<�^��gb�G�A�ܾ�z&U��Z���D�8�dvؚcXc�m�w��b�:�����A;�����o�RH蒁��q �-�b��]b8����:�Qdԋ�.�����!�u�w5/T.>��0��U�t�h��o�5�u3���f�d���
��ր-Q]2F��K����R�w��e	�S���K.B�2g���O[��^���݁G���_�s�~���k�e�g��T6��"Z�PW��+���Ɍ����X\9��aM�b��2�Q����$�S����!���~�L#�)T����DԽr)�h�BV
�<wd��,,��q�A�<�jO��Ӂ��v��D>.ϱ>��"��Ql�52*��^$��'��g�>�r����]'\�9��9�n<������>���Z�xt�c:�(z�G!��(	���L����@v����+j�NyYK�Gw&L3�� ���]���Wb������_!��rR��{��a�3wA��&D��~�[4 �J#���4�#�vX�e�l�y���]!�\s@sSQwA#����Xpx��}YP&p�U��1���Z�d����J�ì��\@�K�+)�DXzƠʈWV5���2]���6��W��?yR<�5V'84t�r�Dqu���n&�_���Nv;��Ir}��k�{��/e�b�%?+����pj7���D]���8�'�m���Q9c���
Ɲ7;��6�v/��G���4ӂ:�1Mu��"�Ɵo�
���Х�>�����s"f(����kLS�Md	X�۔Σo��u�S ��ɨVBJ�JN#T�s>�qny�&�e��sTD=*	-����	s[�c�̛_~Y�Q[cD��:1l~�x��F��{~O���������V;no(P�d~����>������D�� R���f��P�y�K���jC�l��t1�U��n�S�NȖ�%k�#=�P�[B�f0���0%I5��BhA�������L��&c�mM���#ך(�qWM�`��C ��_ �~r!
[��鯸ZE��{���f���3`�M�3{��3�8G�.7J�ޓS2^���{J}c���͔�m��OS�(����Qw'�Y�u7;�JXGi$���:
�jq�!i?~,U���@?��;u�9�2��5G�3^ťL\�Y���܅7$�%e�C�	��%�ek�F��bv�淟�]���Σ-��#�8`T�����)T��lR�d�����D>��/�}}K��rB=��[�d|�r�S ��%�}1��[П	���ɦr����w_�e�G0��0u�4p������*G(�u�<Ss�w,$�V'!��h�Ix�DZi�v��r%��
�J����T��L"Mg_�r^�!h��R��	ךb$0�館x5�3�-�KG�6�90��9���7 <�̘ƕ��sH.r,�Y�:z;i��|�LМn����+�tK��΀<z�'�iD�! ��	� Jx�
�4MN�<�D7��$�(���q�!�� �w����Q,������e�	��M)I�nе�&�j"2/�Os�
b$~}������Eq���YYF��o5�"O�d�g�C��cga5��^ܢ� ��E�!:
���M~_��'
���a����c%(��·�F�8���;	��Ј���.�~w|��aD�1���dy�C����PL�u빁Ƹ���'�R��w�>�����ý6�J�Y`)��Ct�+�\p�~�x��j�M$����s���_d�F�r�~�!��&�f��΄E��]n7rz V;ps~	�>�O�'��O����W&��DEꜗl����)>�l�=pG�zQ,KS/4��"�Cs@OX� `7[e�W'c�A������ {:DN�#v�1�\���5�	��:1f{2�K7Q_�M(5҇.�R��� Sj���	?�9ÂI?~�s�����R+/1�Qڹ�<��F\Wg-4���ݪ�tr$�3�/uk�3ϴ�����)�U|#}�k�K�����HZ��$jS�h
�T�έ�����EG6��O��?��t��	�J��X�w���oU���)��u�S���/tSF(�8�ɉ�L��
G_1��ur
N�5n���w.�_��R�>�7�gIb|���5���`�p>�g�B��;p߳y�pmP�Ngf�n��X��(���&�hq�P�u{J�ڟn]����u-/z�²�"N�-��%�6 �g�֋~�{O�Pau�ވ���ͥ���N��tv��i-�"� |>�q����d�'����?��+1ߎ�v�>������"f����U�R�Q�F�1�D�������k����P/V�q�͸1����'�k��B0���8��g��	�J�؆(�'i��0˝��q�[��y��a#���EPF��d����y�V����C�UD���<0�Q�>��,��R B��8��2n�͘�ɔ<'8E�� U�-U���$!AhE`��d��_t��pF��B�}*��Ӈ��,���۸�E����b�f��[Un��,^�F<H�AY)o%���a�^�{d⁲�%�!d�.�G�V�Om03g6�_�V�=R�0�.yA���d:�K�	T��ǚ ۤ�j����Շ����7�߉�?r�a]Ub|Yy�� �s�"3_�Z�
�Qu=n�ε��k��LTp}M�"�]�f&Ψ����,�I5����ǏЖ!́���E	L �����I#��.�}	�Z�ҝXN��|���we���+���b^T�#yz��I`�qB������ݎ&�>)4���ߧ!�åh'�H�7��S��q�q�����$h~���b�qȢ�/�'�E�p~�j){�0��z� )7E��W��-���[��d�A��T��2����y��bF!x��.\({b�����N��������)��%縱�y!�&��e���Wun*t��Qs4id����(n�g�< �8|M=�5)�/v���d���A X�4q��U�2lƜ���1��`��*{�-�@�T��*��(Oh�b�RA�r2�Z�8�'Ȓ��������W�j��3�p:��^`|ϕc9�}0f��������c�K�/�Af�Ff.���l��9�G'
����@��򌸇󸸨�œw��7�7�<�z�pZB�\γ{PlRV���z�-"�n!:ᰛ�O�w*bS�1~����Y��@�?�:)4�98�eP����������;F�Ƌ��}= �p~׆Pk#|�{`E��Ql��	�f/������ݼ!_C��͈��ڶ�v�v���x��k�G�hv�X3p$ǖ�ߤ� -V�Sx��p����6
"A#����1"���;f�E��A{�}����Q�����1+�s�d#��H���rO蹅�MS��x7��`3u
T��LC]H��A�����o��3�Ux<\ժ�_�B3a�4
�ikX<���#�"��	���Wkd�xf�N��j��k��C�H��o��a�`����2�,Z�n����޺���'�0�)���,��7��&�TW�N����=3!7m��x�%,�@�m鼀n��V4�xX(���u�C���D�bq��ǻ��R�������Q� ������M�.����5�i?�Tఱ�wE[o�J��Q����F��!\FPQ <����u�eˠ��G��^-lCS�¯��+�]E�� ��JA��?̰�Yu�ؘnnR/W�Z�g ��ԟ���Zm/**nb�c�9�n"/f�g}�2<�k�{L��yH���Gq��0U[_/gҵ� $0�%l�K��?��Ǒ��u��j�����2	x��g����إٳ�J+Kn>cB 㑪H #�y�/� `:Ѵ0z2Uݮ��`��[~m�MQq�;�~&�e�� �P�ϘV\V���}]��!��p[{W�>��v�lKB�H�V����~8��s߇��2��G�b�m��G̃g}zǶ7�|}T�$o���ٚ!`�����yp�~��u/ۏv>�Gg�0�М���h:������0`��p���Z|U��/�#OY{�d�w@b6�`�Zֹ�HN,S��v5��`w�QG���R�K���ձ���Ėp����d	�̅[G=�>I0��ɫI	RZ��.��#�؇W�-U:� *ԕDu#M'�?��Ĵ�4�!}�~_>̿���^�MyΌ�&��#�a+�Z�G
��:�n�M.nPv�sa�җ,�W�UC��F���XE��xq �vC{�gX=���eI┆�k��b4|��6�Rb��L3�Y��";��e��d�B�d�)aT�9��-C��>�VI�T�d7�R:��D��X��(�/C���&*+��}��]f6:`����q��R��wB-�P ��*#�v��0�w�5��V�w*�P��T�Ԃ���#��cc*D5�y]�*h����">����yj_�T?u�
���B�#�0F�x��vӿ��ICӚQ�E�=�Ua�z���A�<Y�=Ɲ�k|f�~�"UW���= %���	��Be���@����(�������<D�%Nôr��4�9��v�l8�S�ScX�4�7�l��J{S�
]�Bť9F4����}���P`f2t�'�1j��͟�;E�\;���_��pR[�� L,e����f��h�I�
+�V�w8O�E�m9�i�����{U-��]�Xy��6/M7ˇJ^B��!V�V��y_=z?e$��,z�V"�G�ƣ�3o05�w^��UO����YE�8/k�]�LmAnFET0�M9-8`��*X��@6-������jփ�*��.�H��$S��c=���*�Us�B�p��DǕx-���9|kc��:�4P峟�&ZU�r�}�|&FK��%����x��L��.�Y`J\��� ���8
�{�սPw�s�3���Ar3Pxz��_��nӱ$�ťrLH=��m���M��?|x-���/�,W�Fd��\��d�*�ZZ�B�,��Wd��ί�b���+8~��
�ډ���x��>�i��E�?7�C�kZ�s.�fC~]�D�x���,+�5��4~�DcZw����^�qo�T��ĆQ���5ַ���~3�>w��b���]��.���3�^x!L���@'�e�}�zH�u�D�s��G~�8pPJ7pFu�oBm)1�g䛷a�<��v-��1����Ѥ��Zo��Փ���2
�6S�%�Yw�uO�1f;_�e���21�<�؎��տTs������{��b����i�i5���
���+�tHiO� 9q�km�9�k*��Yo�n������#�D� �uC���zu�&��q���6b�kuذC8{���AOA�5�|�Fe4��ă�<��"i+L�������v%zE&ky��a��[_��?:o���欚t-�ҳ����x!΄�;�:L8x�Wҵn�>}�e�ȫ۱_��c�?��'��D`ɆơGlz�$
���tת�C�`z���������&���׽s-1F?���7�&
�ё������r�Z��[���}X�r1������􊅕-�^�q�˫-K�YK���=B��	Q�[|�F<X��%�Ѱx �l������|J����O��QA�o��z�Wa<!��,]d�IH��Rȉen�����!*���Qz@^��C�C�#0=
�1�w�ܸ�φ������
�zB*�rr�f�|�ґ3;��i}u)3�o���N}�6%93�n�c���ۍ��$��g<��|��{w^�B=0L��O��w(:뫦-�����O�R|iP��3�x�L~��(��iX�s�m:�ۇE���Am�QPi��x��N�@EM%��َ￀%����=���o��T���ܐ�v좍��[�C�"b0��NC�c��6���4�f�i0v��V�������Z~C���Q��`]LK>�����s�Lg�1;�	/�6�S\J��$5��#<���k#�k�	,��yO�Ѵ1$���ϸ�Q��1I3A��%?�u*��o���[� u�{��� d�h뎰��>`�cR�é>�L9��6E�B�*oF�E!�I��4m=-|��y��C�r1�mԶ�D�3<#���ݿP/�'�Wu8����H^pk�����H[I�<l?:��Y��y�^ u���=>����O=�ʔ3՗f\G��(# ���<x����,���1�@��O�s멶��U����d3O!mVo2Ϟ
N�zV:n�ö�l!�kw�d�0,���	�o}L����ښM
H�Z�ܶV��D'Q��AV��0o��W
����Ml
��> F�B��ܑժؤI�.��|Qɉi}��oj	Kf�lVR)�7������gg���Ҝ�AzH�Q����N.��ڦ꘹��t�`�C�?�ۇ��=\K�fk�����yG[��\����/�Eوl�S��+ob�&Dqdk��j�`ʌ����7h,+� )��@-.�nM����^Y�(/B!�0���H$HVo/RW�@S�
���Ų~S��B���?b���ೞ�´z+��:d?_@
J�3���s3Q6sU���\���mؙIޭX��G�o^v����*EvQ�7��8ќ��s�f(�3�۫>� p�R�h��Q<�:o�"N��y>���ƌJ�40>�b��+�X�]�o��$o����I/]bJ���4�d�8�>��x�^ius緕`�M�U�/��<Qr=�[�EG�KQ=ɇ�<���ߣ�=�+���.��.������gY�b�\s������0ܖ�7���1#�"�&��9��P����n����;�P�;�-�����v>;\���5���5���3�ﷹ�a�r�P��Q�>�����Fd��h�M�>=Q�?$�fg�2"L�BD��Wm��C���5H�/\`5޲^W���/O���u�F�$�����tT���fc�mǜ65���r����{\�UCOGZH$�X?/+�48���Ё
��WǷ�e� '�mn���E�N��i��t�?�>!0P-��F�᫟ӑy��T�� I<Pe���ߦ�5(Ҿ}�[W@_�6��d��~#�w�t1+o;L#>����P������!���-��O�:�Y�]G o}��b���(����!*�6��N+�$q�!;�7C�k &�A�śSؒ��H5wu�ڹ���׏_����i�?�Q���:�U��G����@֓-HM NB�ˆp�),e�ھA�\6��!u�I�/3�FGՎ�l���$(^�$�Hms��2ÕB;2�f&��a[���9�#�����M{��ހ�o2�L��Id퉲%�v y �w�#�R��Su���.7H!N���l�� �1�װ��y�� /.1�(�E�S:��nl;*X'��Xmg�����A��Q[j���� ,-ar�*g��@�^�Ef��;��/�/H?8b��"z ~�y���Z`+v���}��Sᬕ/ M�S��+z�k��3]�7g���m���O�Ŭ��h��%��F�MTB��j�;Eso f�Z�(Y�����^6��!�� T;"���q��xp�P�J3��
o8œM����9�˓��J�
������U��N{��A��}~�O��:�7��rb�Օ�k-A6mq*O �Ӭ�_�O�8��aÛ���#�u�����B]�l�������T���p��N&�w]HTFÇ\A@�u�z�6Utk� Wy��\Qpһxz̶>��oZ*�yE����j⭏�zĵ~��rSR�|KT��D��V���Wd`���� ����X �w]BtcC�>��8%%j3I�%��e�����[�A�G�%�]���sR�0n ��ݗh�Y��o�t����F���J���ϰg�=6�g&��o�Q�/d��K��9G�E���z�p���CC�C���X����Jf �����4Ĩ�u���K@%b�yɈ���\�]0�bo��`+e�(��!h(�vL҃CtQ����6X[�C����(�8r�y8��"����Ba�F˹�v{��zp8�[y�u�B̀�G��&��f{�		é�7�o�.ˋ��S���4FX0�\F��x�OeGVJ��'u|�� zW�-�^@�a�EXW���ՇUX1/�eU�R�.�a��iW�K�f(����\�ھ[S��z�˩����:~��eT���HsҚo�$�Ur��ʔ�V��]~~h��_��o'���cwf�K����5�L��̱��G�du~ʺq)be0�mzA5��~�k�ɥ����86E��d���[9����s�ٞb�xەC��k�ȡjO�,G	/=��-o�5-gU3Hq�c��� {�s#�7H?�[Gm*��>9ר�7:���g�ѬWH^��������5�a�>����ҝpbEV�0*ސR��3�4�y��o?�] H2r3����%�͟����&�j�ġ>q�Yy -�iV�gT%�҂��7�襳ޯ�b�8��hhI�
ʖ�>�&F��	JF}�TA�&��J&��	ĦpK�Ư�xQ-��)�̈́gVAV��a��ճb�����egg;��Wx�8�(�߱��PEt��s��b�Æ�����b����D8D7��<W�F�����g+*E�I��[�2^!������	��A6:�p��^�:��f�)']./��6�$QLY�:S97�c�Q+��Ա��*��*�7��OPtB�拾f-�9�tcϱ�� �)F���6�+,D�Ƀ�*K�p�RW�5�qD[���]��Ƥ�2vV���OܴE嵍�!>��tB���.�Mرw/�Js���B������J.��
K���Gj-���D�e��)ݿ�Թ`��Ƶ����!F��\�[`�F:�����E��P���C}���/$��C�)qX�%�`�a�ZvRmu��">�/O�w>���/�L��z�n��_C ϯ�!�U�M',�8�'��J=��{n�7�����4����=+]�]yO�_�:��hf�v���vRze���C��{Tϩ�ǧB�{y+,��&�z�H���9�!��V�9B��t� ��[�M�Xuff�% ����jk!a��7����(��i*a��cs�	'�U}�}n97�im#�Ӈ"�����H��g�،��;������&rY6�_	EO���A���Zv��c+6}'�y����bQAK��>��+sb_�/���k��f��b�R�N#�˘�KGyz�1�4�!���JN�Y�{���e*�mo#�τ���1$��t�RP���u�l���E����6�	R��⧘/d��2Y�4��;�KH�@]�������Xen����a�Hc�
��!�F筎1�?�H�< �&jZ�P#�]�+��Z��UTb����^,7�@َb���H���81��2�A����{��V�R9G-�U�k�v�K���?�l3��|׽��������w"��C���ZsܺKg��>@U�a�$�0ek��!���~�/m�'w��5OF�i)�~ؐ���{�#"K	�����*������TJ�W	�������o- �Ԫ��yU�{+�V�W��D����]�,Z5_��X�ar�$t8�'��2-I��=¸xL&,��YD�$�ZYuL��KLU�,F�o@_�f@؃�!��;�ĵ�~�ʹ�p�0�˂��oh�{�߉Ҩ�B�o(����!�����)�j/�(��XE�Uy��[��e�X��߷�d���4�]�Tm��#���\��2��vZ�O�eJ��rqܞZ�!7u_�EԦ��Q	%���N�ɾ�qK���O�t���蹟�s�s���k_�� EE�P���i�8t��(K?�E��`���O�\������F^#�+G��2�";0lm	���G)�T���su����x`���DbÔ�n��d��]|�r�U���lMQ�n�^��bL���&kE5�	.M6��.2�!��#�͐���c��gF�n��I��@8}��EE�@)��#P��Rͧ}�����O*����l
>�,]4�{�lK���?���|SK�(Z��!�h�\G���JQ�م����1dM����9��+�{H
����[�@d�E���?#<t7��W�p[/��|�\�9�*/zF@�iO�?��G�[�����ψ>�ٶHOAY���dH�	N5��_��s��W��Ep����^�2⇩�F.���!��όlբښf�9�"+���D����=�g�x�U�����8�~��7R�5;��� ��ʫ��Ai����ƖRu�m�� �D]9��(6U��MzR�}��Y�=�Нc�W]a�mz�L�p��Yaƺ��®�ñ"Iʼ��j�7�%*��W��b�p����t��r�FU�W����a���0�+������<�����J�j��3��[�,4L�
c ��Z���<�I^:��v�@����D:C/~@�'һS��T��.p��rB�Z��
rZ�����6��W>'9Ys_j�t�	���9&�i��M2�j$�����}��a{nu��FhTs� _����9N_XI���L�=�'7��,��^�7��/wzb�~���q_K��BiKg����.E�,σ�!Է�ɧ��¬��1�� �A�7�����2�D� :�����G��4�ns���FVΊ���.�oCq���"HP�YJ���AeNA��a�Ϲ�2�4�77{z>/h���D���J�0��v����::w���`��p�{���y,7z)F�K��������7���R�s�lS(]�m�"��3��-z������i=񇟻����x��'������2���!}0$]p�jh�8 m�K��++[�Ā�+#��T���6�� }}�aN��׆�l���4�p��eQb�� ���z����|�=���h�?"{T
���'�E\�5y�Nm�WYy�,��R"�m|8���N�_�<K��|�²z��:�^P�nK�u��UG]�{�Ʃ���U��NzYDBz�ߪ��i���9luu��P�T14֛Z�!���ڒQUp�]Or�'��Gd�V|�?�yn�T�T|�n4����N@i&,^8[G�J�k4����_�sPFt~�?��D]�(��k�t^����K<����X҆�%]�Ԛ7;�P�74s����
Ϋ+�{�K8:c�-�S����<��V���ׅSF���Pޛw����c�x.Kq��<n���/e�ox���A���B�xM��c�`T/�t���k�4.S��_��m���O�ȸ�j�l���)��I0�IOM��{��Z���D<W���}׺��d�^�:����شZ���R�pGRӆR�����ޢ?�^u�IC]��de�I1��Ue��U���φ��t��ݸ���Q��{uH�`�ufC䄀V[�f�}��
v۔}�H�<��qb���gs���W��9o�ڢ� `@�d�h�cь�7������B7t��`��X�C52��<��~ @��5w���/<=�T8���{��OO�ߕ����?�����y*�.�̣Ʌ�M��k�=K�]��Ҁ���|M�D)$�tkx�T��$w4����I��o�^��R+�C�Kٔ6K7>��<���R,�2^�,��>���d%C��qP��#�� �!U^J��6���ӈ6�w�hz%��Q'J�H��,p�B+DAP�Y(��R� �?��Fb*D�w�4N��%�=y���B},O�Mm�3ٛ�����sҿ�(e�y�8��z�`4�?O:ƣ-(>H.�B ��@�:J��N���H���k�y��ۖ<�Q<���R���;�%�%�/�H�s��Z�a3��Kآ�������v��V+U$d��I՝���}Pۭz��d�(�rQ1Θ�+$���6����P�d��~�����4��9r��	S�e�}��ͬ�JW���'P�d���u���v�6e������}bY�퍶7ٍ�=��2�Q�T@%.�@�P���|Z����/�慻|_���zߚSG��sn�\F'��< $k3(��6K��|��+"؞��WUg��p�m��MF@3Z�K��$4�c$Nw���c��'3���lյT�gh�FE�>BB���1-�E,d���n�E�mzЗ4��4���s������Fm�_X��������Е�fG���3����>� ��/��+�%��lb��!{Ǡ$6�?�hc�nLP�Q'�z�W�̦�{$�H�稃�[6����uktS�퉽�)e��b��h{�0����rˋ�������ؐ���qy����"�񓬹;�2Y��N��s�kz��ʋP���ר��el؏n�N�Mʓ�g�O0|�&?���[A}Z�}�|d��j|��!�v�_�n�� :�dZ�6s�ơ�=Ex�%��\��(6��q8�&��M�P/�Q�,���Q;���I��W$�o_Ja���dM��$3�HB�o�M��i��ϼ�����;b�Ć��`�I�r�E�骜Qy���<v�y�j���1�r��Q3&m�a矆���ⱈ���/�!ܘL�׃���G��1�C��et9Hv�r�4���3*���8YH����V��#&�����w���}L��fyS��L��mk�H� l�$�;�k	�I%��r$����AԮ�'�*�_�g���y�VU�K��Ɵ��$ �{��6l�������\�S�B%s�Ӥ��ݙ��b�F6"c����>ը�����Kө��Y��(�pE92T�Cm�l]6=�)5��8�T1Xdt���y�������2�l����q���3hCWB	�om$�.E(.a���7L�*6�v%�׀�#�!�u �h0���d74����x�Ѡ��%3iG�OZ>�R��m{��0�iI	T��j��Ϻ��dhVp�������1�N8è��/D��a��[J���n�0���*���t�U�BL���Z�A���e��ӳ~���Z ���q�y5�!�߶ċ�(J�W�ym�~��]l�^#�\f,<>�sx��.6je�hW���<��h��ʒ�C�r���H0tw=�:�E�7[Ks�nWz��Z"�kh�i3k���ǋ�gr��ʄרTy��қpnX�E�ݘY\H�jM�5z�y����sQ[~�g+S˕�� �o��/�YZ�-�p�Hoqn�\�,~oM�G�9�HV݉��A�ts���L ��2m6�:�k���C�DsC��J�)���'���D�.��c��2rA�,�	(��CЛ���Ay��dR������ۈ!}���@�S���"�����h�H�����C��zU"J��P��
C<�C05����g�,c�f��g8u�j�p%ICڃD �"��#C!�<vf# �Z�y���/��`A��f��Y���TAkh�X�\�F����vɫ;B-���E�؉�9�Tk�.�S���r� O|�B��5�?���+��h�SS��K�<P-�騱��*힝�U樵�u�Ҵ����'�uQ]B���@�n���z���{�냇O�T<�"l�����F�%o6COBw ��@R�p��[�����x~��8䟾0�]�O��O�,�rc�I�^�F����R��P�/`����?��?�^Z�2I>����3|U�ڏ���7Ċ疄B��+o��x��>e��w�u���"Ի�p�*�4��t=�����r�7=�Q�`�	b��y~������*�g6�h+n0�\��-�&��L��u�9��>}@\x�z��م���K��z3����O�R�ar�}k��ɿ�/��聊j�P�;8a��%Ӱ�-.�[N�)2>����`���8�0�x���ߔ���[�H���`@8駎�G��n�o��lUa$ "	7��xcUq�S�f-~T!&[SF� !�O�P@b�(��C[�Ⱦ��'I�"F�]��<��TG�ԗײ�a�6ne��I}��u�h����0?���p4���pu����\�;b�Ls�G���6/q2���D<�X�d�� ��ڑ���*�t-Y�!�6A�[q��m��f�g:GUj��	.D�3����䃸�*bH�b����)��E��F��Q�#�-�ʑ%'�w>��������y�K&deJD��l��DƄ�&pK*���W��5��1ma:pƟ+ *�{�p֟:��(��t��1�
�pN���w~Iu��=<��6��'����?���+���[p;�t��MLm8�x6�b��5F�M���H������UXu4d�^��^�?Gۈ�U�~@�����RYd��a
�I�E��;�t����	j8�I��zy٬���%��LY����zn�X<yY�K�8ؾ�cV:��������D�$/���|��mt���RG	J}#	��.:iޠ��\p^
�*�|�I:�q�#�������7�Qh���v�����9\�Fڜ����`^=�?'���Ѵ⋥6^�EVI��ɢ��(毯���c���"���p�vr���F3�_@ sBa�WBywX-,�����	����7{��'�[k,x��$�XZ�_\�`�)鳊Wx(�of�,�Q�&�7C�pF0���c��JS@��ۭVڽ�Q�Ĝ�ދ��O���:��=f��a�w:�d0�6�[��N:�"D���ٽ_}������[.Rl��V�#߁p �P�6�~+>�N|)����cVzR�� �R�W��=�w�{�]@�%ϙG�m��1y��evרxXC���n����}�Z���.�:r�1��=�(6�8?��¬������/6���7e_��ᰢbW�>��e�,�#�'U����X��r�#�`r���3�k�qE\gt˷(5 ��7	�ڿ&���_��Κ�=I3D�Z�������\  ��Cg��;��7�%�\�(��ӹ����w��
����P�r�Ֆ���2�F]Y����s���Blߓ��lOֻwjµ�K��+E�
��/�����׉n�k&�G�~t� ;%o���m�޲x��^]iA�}Z\VQ���l�I�㬏4��?q��Yk�������E��AZ�ۀ��6� �dD��7��;��kT
	O!��DN�8EOf�����&���vUgl?����ё&k��9�����1{����s��c��F�-0(�=$�Cc�3�*;�v:>����P�1r�)�A�#| d4n��% (z� ���M�-n����T�j^2�r�@E�4���U5�����z�#��a2G�ăo�H�^�����.�w�쇈�Q@����h�����t$!ޢ�`6s�{jy����Կ��;��}�w�Qg�pJU D����x������7�f��HrҿP�cOt����ׯ����t�g!��o��z��Tx�9�<��}<�R9����M�0�u�r��|�� �}����s��0$���F�c�x�#�M�&��e���ۏ�`)��wT�w���*/E���Y7��U����\T�c~��k(���C���#��8
v�W!'c�}F]շ��f]7��R
�� ��Kצf,F�R~ �M�D�:�1�"��'�������=��7�<S�u&���5�=���&��Ě��;��vL5+_ý����s�?XO���@f����:i��fɦ�5�Y��akY��W3�3��1>��n�kA������3P&JV�	�ٛ�>\�x�k��m�O�*�Zڷ90�r�Y`�,h�����3������?z��̐���O(���3���ޘ������4S�It��ٳ�H���Չ4�N��u�^���|�Um
��*3���қ]�kx�R�`�ܶ����	���R�������g��cC��lƱ�T_�Y؝��5l��;��(l:���{8�η �\YpfnjD[�.T��`����A��9T��Q�b�����]Ĵ�7���A��lS�َ��*2˹��Iߖ%��r�l�7ѝgrm7����V������@���t)�'�㭾2��&Y���|E�M���G>�#�>����L��'�	����(@���GB(J�ՖǴ*>�,�NA���1������e�]�.U��~�b���H]F��L���R�8o9��;�b����e�R#]d��Z� �?vA�J�Q��k�M2�w��~'���*
ZG���@ o��oO�f&����Igx��:���	#L�jf�҃��A���g%�?9 �xR��e�Ne�Z˦K�y��2n�s���0]�:|��ņ}�=�o:��ɞ8y�Y'���œ�-@�� S��U� �!ǬObکYN!�ͷ�~t=OGjŨ������񴾟h)
�# 9iZ5���jF�'�9��L��C�ou��٥J	�#�I��Q�<��-�i �tݬ���~g�_�K�3z�t� �Ծ��GN1��v������e}��N�E����X:e�.ȇ��]�$a�
���vC��*t%��O �����Z3/ui+��0�~�0O�����<4F�������c�����k<|�����XϺ�@�<^�e���K��m�\6_t�85p�������E�q�1�T6��
Js�<��8�_jI#̂����4�q�N���-�߳	�iB�k#��X��M ��
��e�Ơ��"0���� ��xR�a���rԽ�y�9�h�a��b�|���b��Y��.O7��-ۣ�ؓr���*��ۃ��j�0[.�S�bX�*z���~�E�m�a$�sfn������F�����ln뉔%�����~ÙmJo���be�H��B��}S�;�!
�I�)Ŧ�`��,���)|b{<�<�K1P�7�"*1k�U�<�y��=�pw�̀��/�9+.#�͇��o=�4�T����W���d��0I9�W��'��&�jz�[}��G�CC�+J��X�2��qæ�n��&�N���
 x�ŏo"�{�S���H^��Rp�ײ�zI�BEC�����^����C�G�B��2�9�o?�g�ކTu��++0
+V(�r:'�P��[SA��;�\gzs�JN�+A��]�<0�ڡ^$Ϡ�ǍT&��#s���7ii�.��Ո��lә��&�WsX.��_C�h~�.H���ھ���d{-^�#q�l�7���:"d
����D�*#��})��q���)4��k/��FxI˖+��H���z���<�����	o/8m��W�B��k��>J�a[�rKí�����2��� ���&�����ERsŒ�����z6�����i�D0=���9�<����U9��� 2�K���W�}�����%��"��y9&² ��F0���=
�y�M�������}��=w��AX��!��HiR3�.0E�Ī�,��B��Ķ����0���.�=�@!�y�s���rdP��q�p�e&\��(֮~o��n��+�������@2�c��?	N���_�S0���|�e��D�g��~n�Y�X���4�)�OT����4��_3-���6C����ef�бb�v���Тa��?b�m�����i`�7L)�Ȩ�4m"��W)�͑ǌ��z�e���&|��A�	�!/2�4:-$��5^#��J�
�AU��Tt�5�G�2QH_�IU"�!�*�����6�W���ƴ�hփ��Pr�%��ja�2��M��)Q���g�V�z���q��3�)'���?Nl��
H�\t�Z��
��P���=dr#�~�:g�=R^Y��l@3�	������oi\�T؝Ag�fMe�4����������!N�D`�S��S����.p�I̢�¼V�Aִ ���J-5/��Z���}�kuv�p�c�ڏ�2��3�,O,;��:@0�����:Q/D�_�ea&c����l�U~:S�i�����ͯ�pz���*��&�B ��T���˟d�g�1���
���|��R;ضU���+0��B7��C�Wu|o�b��Ak��WH%��z
g� Yx�C)�1����V��Um��L�qҘK��������B��x��������!��Zn;i3���ړ�o��5����kn��l@ʒ� �)l�q�<p}����O(���ފѻ���L(Qr�� ��xa��A�Tѻ*��@D,�K]��7w2�؈
� ���[��V��1��7�D�y�%̷X���:��?��?g;�X�`{��|�Z�Y���qaI\jd7� ��� ���Ւw^���6SB����_t`rc^UZp�(ʙx�;䕰֚c���Kl۪Q	�)��3�v^%jy�iP����T7���+/�o^7��R'�UTx��0�>R�a��p��:@Ii�i:%�@��Ԝ2oϿ�:�'�5;��e�nk�Ĳ���Tm�i�K	D��K�<�������l,����?u�-�;w�^ �c=>I*=��x�&�E���7�J�z���x�Gy�lp>�U�q=�ڮWB���Б�;{>lr%��?�����74��LRu;#9�aj��r�^�v��t�e�s��7� ]�v�<�^~d�԰hlV]=��S��wz�2�����
�;�L�1�u�r�+Z���Է�Λ�ؗ}	���:l��jԍ١��P���4�yɮg�Č�T8�㖟��"7H��e��r8
��TdGU3��It6�����P5r�����J�����Il@ ������?�h��(�����J�	��P�p� �F#��s��gR�fA�1id{B�J����Ԛ*�L���Y��%˖Z�n�L{@-�m@5��4
�8���O�fǻ�i}��P�pƫ�݆�ӺT��e%��o�pBY���Z�j�9N!6qR�q�Y��d��-�.��1E��a$�Gӷ='K��ݶ��;4�Z�gz.���M�O�FQ�u`���H��{�W^��~枓��EQa��В�W؀����ᵫRQ��RƄ
�
���
k%��#���	3w<�K�3Tl�C�=qNUhD�ƐF�hT=Q��1�c?��C���!�E��if���kg�6������&�i==u7��o���'VH���:��y,�w(�G�U�|;�f�[$�YggL�L�bM�� ���ίu�o6)��Y*�9��z�U�:(fOU��w2?�S����}�7�Z�PQ���EבN���7Lai#�r�w���9n�S��e]#�Lf����K�y�'"��毠���ĄR 1.X�18�U�����U���}|t�14k��|T�	�$�;�$]�|�܄r��͐�s�^/��<+Ht��=�LP��{x��\��g��Չ��R��{��7�5Mg���j{��ņ�*3}`����֫*�j�ҘE��A�w�L״�Mg��'��0�v��A��@v���F�Z�	ؔ�r�|�b?k�����t9s�R�_c��/w��v����\L
�J����}ƍ����uS:Yͺ	T�r�V���!�CCBMޙhq�6��B^�a�:T������`5�ت��4q����%�������?Xq��y�.�����7�W��;S�'���(�+�hw�߮%2n�*�Ӑ�&ߡ�	��l���Tz�2��>�����'N�n�s�A4/��j"U�C�cÄSr�y&2���W�_0'H��<S�C�!��rţ�yi5J4,�떈v��Xv�h������S�.J?�Y)��c���M�"	����@�Ae-�CX��M�tAxD�c�A"�����#{�脍	z�6�j�Iy�����{jc���I�~Π����t((4�sw�2�q��Ѝ����9�;ͽ����z�D,�Fhx�y���R�����7ŕ�d'Y�_�v��z�D9<?rU"��ۺ�rQ´;Wj��ג'r��
`=�me��՜�鏐��ZK�����G�:����c���&�3Y�?��\���腂W�7��8��ㅔ�q.��ݦA^>�h!ъ�vg���pu�\����-�ƤQ�V�zN�����]Pk"-v��ϛ������eT����&�P�����4;��G��!Կ)5&��)J�m���=����O�_�l'� ���i=�3�
W���1D��5 <��_gm��[*��Z ���L�
֐%F���� �`�-]r�^m����h���Q{APn�������-�����_���������K�φ`�_�Jž4?��cQ'Foѭd�?4�3���7CUr}�&Bn��P��fՀ�{Zl��e�k���ԇ[���X-,�L���l��S~ �������ˑ�b��)b8�w>��ϖ$&�[ x�}�}j���KFP��ْ�n�f#�U�iA�#��2��u}�rЁ�`�[���.�I���|?v��{�_,�����p���ܧ�wq�!����l;�:�Mj�@������/@�XH8�������Е�J8�S���e�\�K�U;�V�Ԡ�K �Jǘf�fѳ�E4ʙ�3�6Ƨ��eR�8�5o�ة���⮂6�h)�J������i�3�\��Ma(!���7�7�l���-�g���eJ�{r��w5
��DB7C\_�p_�O�������@4N��E����i#⌈9�K�f�-8f�P�����M�oE,��aN��'�.�;��0��z(w��$��S�~�a��+E� � Ke6m޵���Jb�p�����M��L���n$6��c��Dr�^������
V��jo_���]\�+��WW��A�/o@�ύ/0U�LY��	��b�;��ɉ���\���U������o7}o��W8����Y�����߷�}t�"�`�KR�7����Q�>z%@�=�(�)��1#ˢ[�oU����-5�����c�7��w��r�����w|0��X+1�綆r܏�ߢ!���{\���ǩB~�ضʙ��#ݓ2��EZ�K5�_�TI7�L����Z�!�������UF;�gI������˺�UV+֚~�WXL��8^��9�my�Ŧ)&_��� D��V4���ȧ�����'7e��S��������~�v�	��1]��D`��ҁY�d���#u�Ⱥzp�ulv
���<s�*�]��_^�P���`�}�h�u��8���&?��M?Z��Y̆=��B�{dv����-�'� ��U^�ſ22���E=]�tD���I��'�	�� ��]��@'�T�Vub�Ւ�� ��J�ù�ĻG;m-�䘥1�E�h
�������;P5���{	t�'�7�؂��,u�A��8�a�\�߹t}�@��&�K*fL^!�X\�p�$��OC����A�0�'���q5�,%<VOȒ|�� ��׊2-�&�bfᯅ_f4�H]���<٘@��0�J��J�hU��81� �ٰ�H�t�<�_%���8�s�!>5*q����U7?�❇Op���d�z}>Ϙ�ɼ�7�cg&��
��
Ӹ&+|�~��u(�
���>5��Crr�.TYRF}+�����m��������з�;���[�YQ���]�ȕhv*����0��'�P�qfTPÉR�0���+�&˂��~%�0#y�{�F�������%�I��&�y n�cH���pG:�O�4i"�#�J7l7�k��
F�T4=E�*�C�J�T�cLQ�p�D�ʨ�&�"��@1��oLNt�Ju����hx	�H��=\��+������͐@FTE�=H��a��xȶ.]uM�x�j��8�!�|V��I^�uj�ʣ05��4�� څ��n���l�h��K�K�'�Q�Bp^�Gx�)���y������h����yo��ܩ�#�H"�yYL������ˈI�GN?K��R0%i���y���8n�>_�F�v�(�a�Î���:�V�q#��(�'}M�xE���$\S3>Ĉ���	�f$9�×��t;��-k�5�w,��䷵jK%�?���ϯ�1y
Η���c�YB��1�3��ټmw�����N_��0�RD�����RO�ʂ�}�e�6S2;�~*��ڡ�2��[�~� ��8�W�9v��i�#B��k�̸0}���	���2�����92�{��S�gv�%7^1�ҭ���q;��0����5z�:x�a/���4�'L�y1MH������A���F��co�ֈ��Ŝ��v��U�lT�;�~�r+�>���Kޗ���4y����v�RqV5�����>�߲�7F�H��EUꂷ�s��7�37� P֩�#��F��i��\�-�H�R$Z���9�ȾI�A3� �u��Ũj���C� ��ѓJ�&Q����E����
�������!&��)��l��H���7I��KP%PoS���{i����͂�[��c�;��%��u/`�>��R��y�)� ����L1��W��31���kx� q��{�/O5? �ƒ��Cu�3��'������Z����xN~�,zֵ�b�o�x��]ҫ�[����v�_s�]G�S����.NH�+!�Z,-�MeT6{��u3��iˀz1�lr��9�˄�XI�-SwW�WO	>��3J̼��Ht��h�36�9���P�,�Ղ�&��@���[�!�[<q�­������*��ALV�ċV��i݌�e��44�G�I�
l��C�,.��Vǖ/_;��Q�s\�кP�眜�@�4��^�+Q���7�C���,�}ܨ����3JZ������9�t�P�d!�A�G�}����׈����Ǒ��,E�Wq)�д�o��ڋN��/U,ޓ?�*6&q��$��1W�pm�N1ؿ��7�
��1]�*pVo6w
�����
���h��y�H7��
M�ɿ5��!��,����Y�n�3ޒ�a5��+�.u�jSX�����_�e������&��f�k���J.��]K�L�'��X�6/B�oݯ�ow���p�=s���ɞ������d�:ب��j3`r\�>�����Ϳ��������3��sxx9+ciy|su
��\�+c���i�~���,
���oP�j���d�0�v}�HGJNZr��������0�C	�	�{8�齶�u�EPyqF��0����>NDF��9��D�E/l!Q0t*�TMc�H�:c�^`uń��یCߺÍn�F r"Nż���g�9j_؜F��kO��D��@�S�r�U%U���L���B}�r��*��X�T��t`:�j�/��Lh�tx�ƺ�澛��#�x(�k>�N���o��b������Ne�z���X���ٳ&EH%4�jm�'�È���(�~���1W�k�k`���s�\o�|͢20~B�عͨ��)Eŋ�5�n-#j��V�%��(5��������xI�d��:�d�
	!�<e�\O�B��*B:!3	����� ���)���sL�D/�c�ZI{��dL[�n����=�Z���+��6*?�H
B#��;�:�2S*�96p|�74WȐ���|L�UV\y�ŵN�{nD�h���=!��1����
��=i6^��C����,j�*:~�0�a6��H޵)��u�P&ג� �^��Q�v�"�{��7�Y����!�!BB������>�ͤ/G!<m^����ԧD�f�(�%�d�r�xBSٕ�H�5ފrx����t���^l֡���!� �£��jd��<��}��P���$�]����ж���5�3��u�|�D�s�c���薘r�j	��d�|{*��߿�K��Q�%��v��6��^�L�w�FM�<��t}��Zb4W}d2`�/� /�] w��~:�=R�7^��_��Ԙ.B�����ɟ/�F�<k���9��ؼ {L$6Nș�tp�:�����қ���[j<�A����9I�O�i78����j��sq�=�+!�-�=�B4jrj*+�U���`�	�K-�NV�Fj*���e���`���)��NYf�貅�d:�B)"���:A�2 i���4?ҭ#�Oi�)�`ؿ��=�����la�]�5�+~Y14˨ W,�Z�P�Q�Wn�hE���v��6�̊tc����M���_m7L�C4c^��_��a�5��M��Ř^����6����(��x7�{R]�n^$M%��/�bR;p1�b��w*�Ȗ)�w?�J߭�vQc_r2�a���Nm��Jt���oj�E�d�`j|�[�	I�#��K�*�9�N�]U�C�h�x��&O B<��˜DH7���
�^"�Q� ��<��A�RRM�:��-�R�
�t��Ռ�����=��f���%�>qB��j[�'�[�/��̵��!�B�Q����w.΍��u��$r��db�8�Ħ�S��������LC�5�;+{����X�j!�1�I,t4&*7��	[�~�;�6����`��Mg�U:����1Ĺ����r�]������-<�k)��S����2���Rx�5Kgt�)4���ϧ4�	���9��
Z��e�4Ƞ����;5�j}�����d��:��2+w��,=��(ߕ��F�T8F
�]�
�I�V��l�F�d�ٜ7붚�:�����r%��e�������cbzAU�1�2�ZT�W�]{�G?����A�տ�B?[��d���*�UNg�k�ƻ&{��	��L����c�}ݦ���/��
�D��������q�y�jY;�xyS�r��߉�2e.��	�T8~yQ$N��{��ԓ_����ޜc
�s��R�n�qWN�+HxbXr[fUD29/R�pb%��|�F�ʛT	������|T�KU�\�d^E���%��7�.r'j�˪HR�����F��|�`�K�����3�0��tS���!��oc̕B�d+����XYЬ����[Ӷ�d�� c��q��a�es@3�m[��=����/3+if�#�I��ig�B7}�F�3U�LW�OЕ
�h�M�#�I\��w3�,H�����������%� ?dJ^�'(��l'��'ܳ��$~K%��ps����d����Ẅ́>��d���x";��ߠ6�P�R�L��,��&��^�57.::���v9���+��^��#tKqb�퍹�$����ZC��IR��-�Č��Ȇo�O��R� +�K�����T|F��y�}��q@��j� <7��ÛO簢�۝[�)ey�M��v��
@=!����ә(�3��]�C��r�pw�7gp��l�[f.V�NK�K' ��6�{���1�y���7i�f�j�7(���_/�
�aJ���*�N���a<���i��?����'f6�&9w��L� hk�St��Vm.�H��k��[�ײ/���u�:��ř2�������N�`#�ʼ�d@M'^��̎�e��&��0G����Q���FpᥧGi{ԂA�1�����7��`�%ᆍ�ȇ'DI����T�#���-\�g�8TJ��Aߤ<�)O�4*{lY�NX��.
�Ȫ���M\��[��klLxEEo����]:�+�IfL9t��e��Qc��E��3�ʉޟ��_[�J����򂟇�-�ڮBX���Q9����V��q{".u���[/��I�$�z�����w�vޏ|�-�j��#�n��Ig��3?�b�x���_y��8ךN��uP�&4u�ڈ���Oz�R��A���^�N��hq�5��b`�98ؑT��m1-G^e)��5��������&蘇�#�?'�+Ư��\��D�T���^�~�l#z,P��wW3|���RH�wJ���c]q���7��X�MTE�d9���_�>A�j���)��n��"8ww�ۊn��g�F�R���rf'Ϝ�<)[s��A���Z)�:���߾6хe��x �&���Y��ui���<4�J�N�qnڊ.a���� �P�h�w h�ȕ�&9O���f�Un�lF�c�w~��n�&Qyzdy2��fǰ
e��h��I:�S����$W��j�kF�����X�%z�Q��՝1`Li��=2�1Z����e�y{��V��|t+���-Q���X9N2j!P��[�uӸ�)���_��P��m|����z������h�+���?���&6w��t�fO�1.h�'�������	4�P��eq]^�4ȼ`�k��	��ū��}� �󩬙�ұ�в9��K�\�:<+��w��i���52��]���.�`�&LeZ'6��\��/�[�{��IB�进�y�>�[�s���(p������;Q��bf�8'}h���ZjG8�9�{<HHT�q9�ɟ��p��/AR�L����}�%����nW��<�b�O���Eܦ��~ 6�Vk�E an�G� �u�Z��t�KW!�}f^)>f�qH����Vɩ�ҋ�B�1bd�R���9^\��C
�W68�bǛP�ͻ?N����w�H����ɲ�m���x��2��OD]r�Re~�R2r|$xك���)���e��UDhU�+F����l���Ag�iOB�f 3�9������`;ßc�2�p��7�� �w��2�>Q�|�C�O��G���O{�z�:��p\h�}��,Ѥ�MݞJ�g6"�H,/���E�'����_j-�mX��m ec5rI̗��{����lmf����$���B�x9B9�]��e�L1��Oq��5ҹJuc%�D�'qY����.�z�g{���7��V,<u��Ҟ��xY ɏڒ���s
�=3q�����E�P�Y��}Q�aǽv�tljKjؔ������+��L�%B���B�U�H��6�bvM)6�hƝ���e!Cc-����Ɋ��$����C��>H���i��οmD�HV&c;�{NV��՚�[�*�>)�}GHmv�}M�����-|>�.�#A�,e��LTWEae�(�{�a�w�.���W�ulZUM��p�#8pRg.ocܸ��])���ْg~���P)0���NUioʇ3�M'D��4}�R�&�mс�t�v���阍�5+L�m���md�{/ �ISZ���z֖-��~��Ou0x��k4}�[�E��9�¨���T���'/�|�2������H�L~ev��u��l��5�`���!A�Z��� ���~��C�4I��m�E�xQ\����_t/Hr(�n���:u6���
lV��c�^����g��:���Q��8�O{d���j�z<�iT�Wa��/e��Yu}%H��;.�l���_~,%���(6�US
�9�m��W�}YfY�֢�@0=��=�9�W>mM�5�
�)ܟX`��`� ��	d;[d)2[6�	x�Y�����Ւ��k�牎��WNWX�� ���QI�$i%�S��X�Q�Y1t�l� ��Q�f�fi.�]���H��j���,�4�ګ ��3�5�e�Ҵ�e�X���R�k�t�wN^\h鲓��I �ɎJ;M�z��Jp��$��":q+��
)���U�1Sr�!~��0��#��}��Z����SI2'2�}�,Kdk�[�ލR@��JBo�zQ�,l^vt��*�A�]�{p��8���r�@�E��Z�m�<gG\��v�ԑ�ȣ���;O�65+{�w ��܌I���q��.Drš��%E��v'�'Ϟ�Μ�h&��F���Y���*��8��p�Eū�puR� ����^I��5��r���#3����!K��������T�l� �%E��Qet�H۰��q��*�9�l&;'�]z��7r��尫����C%X��O]r�&	�+�6���T���\>�$�����0�O9dK0�0ݴ�:��.�����my��6�O���!;Xc���������]P$1��c������3�P����
��=t��Ît�)��d-]5x<z=%���P�T��!��v�V<HL��oŁ�����4��]U�y�G��w
���-�I�گ����R��b��#�"wF��3��^��	��&MεvЮ �R ���8�G�|�T�|��h�i��rP|�^����m���t��|e�hjO�9<�
/�6#zj���7I�M�H��� �f>�S���k�%{�I�A"�,Sv�}��0Ƃܐ�R1Se�H��c��L��=y�:��\��S�>8�)a239��J�\���Z{���<��	_��*ۯ��/}kw�C@�%2��J�"�Hҝ�hEod1�+f�HiP��\R�8�[)���5�M'�wU�J�ʋ�"���7���.�G51ҩ�)j﹂Y��$��V��t�y�>(ƈD�8�K���Fw�Mo��L�h�/���{�|�
��gӧU�f͌���$`o����c� ������K������?C�-�����Fr�g4�>����I�Z]Y��l\�p�:'Ođl���rY�k�t��~V�֪�DN�QX��'A��T&�L�>�uCSU�=��.6jJ�S�b�����i(��,��5��P!�����G��]��9�I6�3��SU#m�V�W��p}j���Jϭ7,x�\�~�HOS>O�����J|���e8��H����/Q����j�cȧ���N���.w�c�����+v}�[ܴ�H�f�%�8������=��j��G�ow���j5����dv| &TRn�"���@E�f�ӵ��(#��|٥��;&���K�a���X���ll���eq�G��~��y,�1�7o�����[��P���9���m!P�Z.�ƭ����Y�?c�!�-���hh|��<��IkE$}��1t���Y�(��bUT��)F����j`��H��y4��Վ(�Pz�Aw��L)��y!����[�H��c�*��'�;%0��@���>��,�7�/,���?j1�:�Ia������$4%��4a�� �nPջ�2��5n��VYz�T��`DhNŶ�-� ���UA���|�c���TL��Ac�P�e����#�����Dz� :���'�ﱵ������kL��ϣ�cYTΔt	.*D6����N�5�Hw:�������q�-�l�񬘞�;���K��y/���eL�I���HHӋ<�_R��;��B���p���n���^`��ɕjʔ�l`t�ƾC�� �ꠧ0��o��V�5����	8�q���j�C�51��9xS���0��.�v8�${�.������G�^[s�J��Qsc�}�n8�.�:��5��٘�j��!f�:�N���Q���>9����i7K,�eR�,� c� �:��������-��6��(�t����f����̩�H	>�=ny� ���47g�'�*a�$�W�ޛ�����S�.�o=��c}S�jr;��0<����g�n_�QC��e���Y��4��v� ���q����cБ2�nv?j 
�t�DS#�?!��.'�,�����V��$Z�ܐ��(uF+KY~��T���j cSI)������ ����a,(�Pp9�!~� &����� �H	:��+�i�XQ�Ns���4n}����1)U���#y��ޅ0ե�����r��֔�Nٌ�����ww�E�9`U��I�{K ���oO���C*����������ދ�%��"��B�=R�U_�6J���p�M���cFX j<�ϭ�D1�lE�07�M`5�3�;z+)(tN+�$��~�Z:,A骧���e���z��B�X�Dso����pBU��Di����M)�!��=0�rAҜ�z(�riú�&�UP����*����� I[���?D��>S���39��"�d�-}pfoDc]~�%�L��֐�aI��TQC��-I&�6q*� ������s7u7c��۸]:�$=˧��dd��V����x�f��`RNJ�%�4yS��l�>�mJ�Eb��V�7�CuMT�=��cEoY9ok'_C_A������x�{g��.,:OD#�4 3-�l��n�����/P�f��
W	|{}:���a`:G[Aa0G'��p�[/�Ê�e�y�ԚyA.�@��^�֭���ٞ�k�_I�Y+Nշ�Xt�	��q�ˆ������~��Ic����]�:CˮA]�+:���C[��r8�[�T�8'�-�$}���d�fKa���7�`6��M��F��xa7B��;:T�S	(����B����$O
F�'��\-��IHsG�O��qv�d�bZT�t�~G*A�>?0U���y��V��ĹW�$pY�M���|��:k�e}(yHGa�d>9��I���	u�Hu�`���^��Z�2�*���8���8ӗO�ܥ���.�.�Q��B�v^�ͷq�Yk~_�VƠ�ͼ�!�.P%9�$���'�H�b@@��4�QzJ5��� Ps+�Z��-C�C��`b�Y�y�����u%t;��&�S��`FKA'�,*h#����Sl��I�+]��4N��  ��s�Yƺ3H�*L1��*���Tt���"	}���A��p�s������5��أP�ٶ�N���a�����wg��;_�Do�Όq̍��uԡoXZ�E�v;�E<�HB-!���#�Iˈ�{�ArZ��f� n���b�\u������>��p�9>n��l����|�
�[��e� ��qzU��_�e����z���*1M���������ѹ=��-�[!T�KY������r��}��8:��4�a�[��ltB��a_<+��V�U���dl�E��@�C2��	o�aK�}��Jx}�Mh=~Og�w�!}F��K���{o�����8��~C���a7� `�3�c�k3�b�Y�IC��֣i[�x�Fn�i�-��5	'.�0�����۳�4���k�f�n�
JLq9s.$c��0=�"���Պ�G5B9.ƬX��S/�/w��a_���H��C@v�F�S/_��ҽD
L_-[.r��A��d���.?�s�����1�e� 26������-��u,��풰�fH�Yh̵�>,�/�O�(&CH�s�Vo��2&�n&JC���0)g�����2�&�6�B���^�8��R,�� �U�YQH�N��R��]����o8:#J�!��L�a�ǡ���G{	0v,��Ȉ��@ۺ�
(�t{��k�}Eꠟ ���Q�z�)��G�X�_�G�-��vAu��*�?���Q�l�L p�@�Q^�W�#� �?�GNj��Ć.��ޠ��$*�HT6�MJ����u������IA�B���x�@�A*6���^Yn+��F\����������GCϷ�?5&?��B�RS(2�r8���E�>�ֳ������E}U f�^��I���9K�i5NuJ`GcV4��x���=ga����g��s83j��57)u��Y�B#�?����Q ����\�Ϥ%�PϨf�E������ͪ8����A*@��� ��Ϋ��i�S��/6�3"�YOF$C���.S+J�~ �oߞ��K����-sؽֵ�-mv!!�ys�󖔃E����Q�x�z��ّ�=���t)K�Ԣ���V��i�e��K�s~B0�T��g��^�``��k�V�צ�"
G�ۄW�,����~灔Ѱ�r_z�4���v�R�3?`�q��H|B1�����aH7	�*�ۤ7���5t]�� gw�������t�C�;�Y�39a�j�AW��0ά������ܔ��Vǯ��*�!*���O�#*�T#����J"E�#19,vy����Jۉ���u�PKӆ�6�]�������OM���b�c*���@
NZ�`b������H�/�ٌ)������Aa����&�����R�|ve��LnK�s�3yN��&�B�ҌU���ŧ��ynO{���t����S6�4���0p�.b/z��@.VX����g1+�)�_=#w[g�p�[ZȚ�凐��Ut@ȳ��Pe_���]���H����Bn�.Ү��RK��~ou��3��D��1w>޼�+XH��t�#I &r�A�b71ҭ���=���n����լd.x��E�JS�ڻ ��xڇ���d����.��b�˞��
���PA�����Ee8T#%��l��͠"G�/��ݰ�@{��Gt_��(<T�e>�s~�k��}�{��!��Ūo���4Ci&��Z�nh)��zi�f��P�|�u����¢�V�^1�Ɗ�=�a8�p�,��<���y��U�����(�`/�4�f4&K޳O��e��?AE0�Z!�E�'�!���L�5�q��{7 &�Z�,�9��0RPU���|��F�;&����}���v�f��C*n{��_+wƙ��|���HVU&�k�o+V����ۀ�Գ�����d��f���X"S������v��Pvr��D�iu	] �L�fP'��s!��{D�@��qmB*��� �Zk|f�q��\Kߨ��`Wl4�b"�VG��̒	�������ů8�C��"%mJ�W�{"{�]]2t�<p�-c�?��YV��Q�ժ-��\��W���vaZ(漅C��b�)3�P :�;2k�q��%��ɟ�^�H�b4jk^ಊ��*�ˍ=I�nh۬B�*����%R����1!t\E*�F��m�D
��������E��q�������1�L���"�����Ө�u��,y�˳W��o�3T{h����m�L���O��y���3���p���	��?�Ix�`�w?Ty�Ӈ%�Q�}Yª�Z�ܦ�5�?6j�t���N"w�D%ex;N��|N`_WKG�J?�D;X�WF��|\�6��d<w�&aD����%`���_�߅Z�#�;�E��P���A'̍Hz���lʵ��
�t CI�ǸlW"=�Ofk�'�p:��K`�P��A��b'��*CQ�
��h���;���[qlV��x�qx�<c^>m�Sm���[Ń&��ῌ�'��Lu��Dd'�1 ���
ԭ��é����ShfDl�	�c{�+�/b�-��t��ң��$�Q4<'-�&:�m��E(�&î"Kg �1"&o�+��ø�_���F��l�����@�u��P'`�H.�͜����e�O�,�v>�r�6��޴U�?��c=�
��V�e�Pz�q�R������7�x�/��_�K�>ˋ��=�?!'����f��lLY���ЙOLN�z��J��njs%�ay/�SO�rq;?�h&�ӧ�w���ËQCȎ}<|.]
�&Vnds���bb<��}L|k�,�q��`����C�m�!����kq�K_���6�X6@�԰�ƚ���������Yd7�λ"���`7<>!"�V��>R��/�&4q9�����z۫�W���H������xw�5;�k1˾�J�G���'��H9����ǃ�s�;����<V%��7�6�ķ+���'7_e:5)�|3�:i3�0<ܪ[��*����{ѥ��ɴ=�/���pP���NȲ�E��a��T�����hd;Y����e�e�d��f+�5�ژA�E�O���\t�8*���,�r#$@�3� '�-D)C�JO�+��<�5pa���}{7�X ��q/_���ȳ0.qȻ<���J�з�߁��&n7�}sQ9X;ͷKO��*�eZ�*���@�I�>��fG�빹rU}����z�Կ-|�Yh��:0�i��8����aM@U�)j��;�y
���Y�C�ôQLQ�aS�\��LK(⋇h��I��s�(��Լ&�JN1��><,Nq}4����,P^�P~L��}ЋU��ʪ����l�Lx��øuܜ����2��r�Bu'h?��E�i-�����-��v���J�+V��\S�5?��?V)�E�:w�����]�&ˉnŎQy6T�)�Pˉ� �PSg_��2��o��b�ǣ+�ÞD���Z}%/s@E�C�R�e�[�,$����b����D�*�4���r/��J���yk��UZ%Bj�1�p��jh(�`��A5\�M�EZ�<rr��E�V~3���a*Nלy/�
�TYf�A�!v� �����p��K
��#���x��и��s��4W�����+����R̎o�W>oP�PtZ���R,��3��T�QQhBab�
Ḩf�~9�l�n�A�g�@�&�'�׋�̐�no�p�K�0։EWY ���B�E���5�#C�E;0���Cmѣ,�Ƨ#���F��).�u�Ü~2m�N3֖{H�߻ ��ȡ�`ڀ��ʹoTɼ��V�)�]�[[� ��3h�uP��Bv�D&�J_<�r�?E�pF&�%��KE��Hꔿ�8�g6,
P�V��O�(�v��P�/�~P��Mɟ����^[k���!���D�Mt�+�y��+�u��\[��[�?�o���L�>�9��5�;U���z�*{D�9������sQp�qQzLa�5����_i����H\�2���kr�u��R�Û�{ �t��4d	n�f��O^�ܗ���)q��R�I��S�Y��QXS�+y�e�Z]˃�	��:⏎�ɓ*{1�Z{N�X�-E6��j�w�+���k��2!�C�[�N�ORls�9����A���7ĳ��;!�\ƃ{c0v��4h:�k_�_E\D��t���,��Y��`w~�V5z�{�m�&]�4R��Qu!�ŶK����2��}�@��`�6�]1L�s�r���8�*��J�7"�c�����o�Q/�ҽ
ϵ<��s�La����|�K-R-fW?���w��G���এ��Q�A��� � ڄ� ��[�=Ly��&��J������<�a~̉�!1�����t��[KEǢ��,��Hf~3�eM-|i����-@��s�8u��2��n���D}_�B��58���C�}�d�k.�SN�h������0%β��	�j�[h��I��,{|��������k~��H`�t�;g���x���S{���Ɉ�X�@�J'���= �n9S�ؓ焪J�sx�x�Q�5.�D 9E��d�|{b"��崏�G��xel��P(�v������l�`���^L�η�>��;�!�r1a�g�i����hd*Z�����s�OIG�-��'�lG|qhU��r>����ܥ: ,2cW��UTt/A%�9���'����1��n�1@�R��7��*��A&���Ɲv'p5
��/̜�*�/�h����*6�ekK�+Oj�.�(Đ'(4ѹ��Ĺj�xx�أ�Ι]�.�g��ۓ�L�|�Z�('�${�m:���|mn8��ϥ��(���m5��T�t��ͪ��E��Yt���1��`�U�/!H���@w�;7��O�cR�hq:���=DmL5k*���8� �J�sN�6Rc<]��	��}��dn�P��InN�đő�͕���/y^�&�B�U7w�3 �Z���I�Y&�M��3�WHM��*�� ��>������ !�!��"!���ZM�Y�Ǆs7= 
�Ɇ�����GV�Q���<�!�����6-T�l]�r�!鎆k������:�焴��N�-Ưz�v83��k�P�7	Ì8��n��x�E�I��/+�t�DM��J�siH����.�M�Px~Ŭ���X�hʜ�̴����:I�0��)DL���ֲ\�@��	g�s�t+}�� V�oF椓(�'���pE���E�+[�p�r�EŜ�l�+��#\т|��:w�T���b"�<qO!n8
�e�F��8�lj'neڜ���r�Mb3o���Q��ˍ��?�sl�8�7����B�?},�/=s�Ҝ�k�A3��<��zT�٨��[��ʝ���6A��7���0ˁ��o����ꚁSz��yt�v�2!�JJ����t]Z�O�DC�����7�1�Z��K�5�< ��Ҡ�xw^�vP�j�;�3)��?�r��>��/7�6Y�j �% OA���&+&�rqV�8��O�=��f�l8	`�Gx���̌7U[q3��1�Mtz�BŁ%Y݊�^�1��*�\�n�k1�B��Ac���
/��[���Nʤ�����O�Q�����󕇔\�J)H�����m�E�Z
�ya�:˙50�c|��3os*Fey�{�edO4ݳ ��v�_�e���!b�<���'����
�7�\gsW��s2c��>Yv�XN:��}n���c���G���hk��sr:�Ͼ_h���
j8B��I��O��&�
�k|;$�~yVZltk���D��WI��<3	�n������2��O^��Q��}c�"�L�ޫ.6H�y�ܘ#{j�"M9��Ղ��z�Lܜ���3���{�8=h=1����$s}�*�|��Hw[/?~,�_��b�d�:�&Lc�
������#f�h�� �@��K�s|�]�̺������SX�0y����brC�&��V�.Q�K���7X���z��lO!�Asݠ�&"�
>�TUp�C�W"�
1�!:v>=B��lꇈ�$�����	A����I��CP�4�����)�Җ�Z,4̀h�3W噕Z3u��ʇ#+lH��zk͌�U�")?����L���y��`[��;�_`w�78u4An?fi-kxr�U��_���2>")�m#��]��*�Ԣ,+�����u�9���e�c��$���~�a�z&��Q &6U	�%���V�!mjN���v �1�X�Ckp:d�ҧ�$nW��w�+���Id:�o���ہ��5�z�]�7s�ԤcL~[e*1[1JT�����������WL
�@��K)��(^
^�f�|R�x���Kx3o�� %�8ġ؇�f�%�����p��'����['�c���8
@o�O���qI�����ߒ�R������,��b�R����tcj"�c�4t�Jϧ>���]Z��������E���u٭�W�t�I�y|��e����oC�s�pƁB�>�قpJ���w��=s*�׌�ͦ��/��Ϫy�p}�1ʛrl^*�?H�fQO)����s��_���Ҕ��[�]��-U�%Y��$�ZɎݐT��R���o�-1/Į�se��A��cSQm�y�k[��`r<��p�6���"���uVs"μ|�����J�q�eT�x�v��̺�
���rΎ��N��?��i{���*��o,¤H"�5��O��U�(~�c��#讅O�}����Ă��^��N�r��7+�ޘ����#P��J���A/�V:g\�Hb}�ͅ�z��oć*��zw���];�b!r�����.{A�~�.�I���w⌴�a�:�,G��/H
B��.�p�[m��a������r��
Պ�φ2_�~���l�J�DS�L󮊫��4H�[y
|��@G����؂�y��ɿn.׳�>����	+u>�ʁOe�/N &��2��zG�-�M�?�Z�X���A�m���g�_O@�F����Y���D���]����=���v(#���Y�*'(+���)�<�ꀭ�L�R#@$T�%}��<�N����7�%x�����I�AFg�38�+6G��t��*C&t��1��B�����X�ܸ��WQPu榭|)x�>��t)��v�}���i�Cv/߳���Va�G1�����$�����k�1��Ņ���/�1����[��N�̎l���ٛD�C˴V↌�(l��b���m����C�(�Ȑ�E��k���@ѧ𔀱������줾��Y�zj�����45�*6��odhִ/r/�p�{ni!e��ܪ䟢m �.W}�<�[��;���Qī@��I,&`��z���{�B0��4.��֕�$hOg�����?]���'c�4�u$s0��yb�7e2�6��Ie���X�X�����U/�0���ht��!��4C�	�B��ta*L�yn��|T ɚ/��Er~���6Iz&"���ߴi�Q��R\� b�"���ZQ�l��I�B�t�w���(��V�|��?'06
�<� ��~]�z����?��	�8	��yd��,�6й�����};2�t0�0����9�,5�;9�*�E ����Ĳ�|��Q�ḁBp�@�B^Ǩ5^B4 8��55z��0�F.N[di��~i�.|�n�U���k (t�H�Y6�p*����Y�vK��1Т���2Oe����i���Ch�5!����\�G�0�P��2��<B*|K��y$7����u4���H�Y�����i�kY������k���/�̨
�uV�c�k0�v�>��ŘWv=@��O��ϙ&x�mϋEm=��<\e�O3�+�<[��69�Z�f������e��}��
=�:��>M?�j�h�9=c?�]�� ^�`��I��jvz�s�t��Y%�)��C�x�v�R�����ť�vfS5�C�$V�B��6��r�Hw���M��:IT�-��#��o9J@q���
k��t�8M�g���!��h�=�@���f��rq�F`I*c�]�OT����2f�H���N:>�$h9Ҝ|G�`��")d�2Z��2B4���
��8�����Du^d����bA�iBk�-����iT�m0O�����p��v�솰�-�?v�6�Q�@���5cA��]��@$aYv"�&�{j:q�m߿� �aͅ�$�Lu�}��Ӭw6��.#~�{;��G����RX(2�@P�.Ps$»N8�A�Z&C:,��7u��S>H��Wy?f�i�Z͇Ľ7��	�b��Q<t�'�����}$���h�( W�z�U������ož�!ʠT��4���5W�U�u�5.x�G��-��⊶�߃#n�L8j��>�C���CLz��M$�*��c%��CCX�"�*+�놗\J��Y�Lh��©̗ز��C�sOy�,0���}$2>�qe��;����d'���%Ѿt	�;���DN�6C��CWA�B $5k������y�=��fEſe�:dQ���L�b)@��D��%?�\�W!p�g�����6�������e9��j��o!�:�Zw/���Q��_N]����'����쒌p��uN_�wΑP�c���5�F��z��J#��!]=
).�Y�Q �m�����~Խ�~Y/裇n��/��:�g�>�C''[�n�~:EZ���)���xR4�b.���b0��v��f�9>����+���
��bȁ鸑Oi�Z��B/#��Ћ|��׾�+���Q���A��,=zN�p�kA���1s���9���	����	�-�u�|��%�4<��K�`�F�Q��Ÿ��x ܢ<u�������NZ�YD�	��v�c�!�nCF4���(��J*�����u�&�D��[G~Z�S���R�6L�H�-�&Ŝ�2�B�i��aT�z0�8h|��t��h�D@9�yh�~3�[�<V'8)�� 4��o�)lF#^y,�I&���M��ѕqo�q1N�h��~�(�$e�$�k0<��6�˲��&�A�a���\f��|�ɀ�!,/Mܿ2�IF?!"ຣ��9�vω��H5��-����
g��ԽLx�$Jw3@d�%3��A����8�#���\<��aVZx<�Y�e}�p���+R'ƫ�h��ä=��|M���r�t�_����^�2���7��z��%zk��y�g��g%y�{@�͕��R��}�Č�v���u��<�Q�Q��3ث� �߳uʚ�+5���K���/�:7����$��7��$s�w6�<���~�dW��3��z����Ø�i��4��մOu��\�b��zL~�Qy^-��h��،��0���s��a�}&��@ ͈�g��
L|��,C_�P����RIc2E���5d�E����m-;
\�K]q)ƚ�c�"O���܄7dN��,��Gh����"_��f��>�k�U�z@��Z�]G�n=�ԩ�����>\��+q~3QR��1�e2TTT+%�6%\×�.6�IK54�j�vڐ�eS�	,�'�Y�~���`��S+���?�
�>3)|�Ld�v.7�����f���"�9c >�(��v^�?�* c���n��3�FQv��l�)��+�X������/ex$�k7$��5����:��3��wt�y��؄#7�7.o��?˂X&��q�%��j��砆�v�돛��h��6FU�h�k/3"����:�hwĈ3�i�]3��0����^��r
bĖN��0�3x.����Ϥ�����'(H�+}}�b+D*jnJAN���9�I�:9�o�1���7�(������Y�w���U�Y1[#�7�΅�-v���$��SI�\��r^�>���lh��SOn;�d�a_�B�FWm�я�d(a�6[�J��ȥr:L����Yn���(�P�1tńNv��,۱�V�wj����9�����|ij�l��R� t�Gw��-�Ó�v�B}���bBW�-w~�fY"���t*!w��ʳ��%��0O9�/���
���e��t\�0L9���gKy$�I��/�ed��2��&Y4Vs��w=��4L{�w�b?��� �Gp�$�%�T��_P��(�`��92��c�2�}w�˳��� n����  
~�Y� ���傤T�7�s�1ڴ��},�-�� zrD�9���Z��r�FP������f݄��^5��=_�X��<����z�� '����k�ĭ�*ׂ:� |]��0O�|��P�6cJ�W��iw�f��y|��7'�\!,9�r�#ֵT�m�~�� m8=�o�\��0�T�wĶ�"�`�%g�Н%�1	�Ԯ��4��=�n@�=%�R�<u�`s�5;��B�kq�$�"<|"E�%z��~g� R���.��.a��svXfz������8fv����s��Z�SD�ւ
�h �����[���]�,�I�.�y�4�J0*��A��9U��������i-`�S���#;i6��7�y���z1�Q���waw�5|c�lb�%��}yP@�&o���9>C^��-p;d�4�@gUYjy�`�u߲�Qby^Q��}{��`v$���X*@�m�h����wS���X�{l�m�����뻡�HG	���;���d>��jXo��Zo��wf�1;q@s[��,3�c��v��M���=1x���uu��(KZܕ/��3��� ��eQw]央F�
��uv;%�Ɖ�ȍ,��lD�d���?!��h���W����ư�u��e�<����e��c�=p�a�Y���W���=pf�(�L[��a=k�61~���O�-
+�y��&Z�p��鎹#8g���U�������-�q�~�珢��o	�Eӹ�C��#���kVs�Rs��es^��CO��ћJ���V Z�6�8��i�q����͇��f)��x�ȷ>o�9/��r�>)Y���sRc�}9�%'?mJ����P�Bqe��'Q?z����-��*sze�ɸnқ���|�C����nr� ��I?� zP���#�5w��jiW����`���Czi:	lV���!��>�rp�ӓjcmtF4�:��$D���2f��P�'��Dx���$�d�>1��ҥ#�m�(��U�����qı!��Z�ߙ�J�{!셄ˮ3Ea�0��ƳNl�>8��3�R<K�{	4�qb�l�tI���e���X5��)2���B���7a���4]i��NY�I_ ��Mz�,N|��U�(��PrCs�JR�e��ϣ2�Nfn�p��!O��br���2�F������bI�]Uh�Z��*R�L�F"���ik�,��i�U8�<�a����Q��XQ������P�0�ىi��$���_��-t5��t�wn��Hr�5Ro�y���$�&���x��l�LW�6˲�h���2�Z<���@�m��D�������cw[W��&���R�]׋p���H����E���qS"~��t0舳�D�|��3�u���
+:du�a��gc���*hc��
�s�pk�}cꞃ��x���3�5�����nelbd5��y����QE�FZh���ǰ'���KV
�v}gr����66�Yb�Y���Ӑ�k����ζ�dj<i�OV��eQٵx��"aEG>~"��hu�� �����|;�E���V7�jI���@�������e�jr�n�+�04A[�P
r�l�����H��{�Um�W��Λ�x�[��Β.J���A��-W�q���E�WjsA�.�7�躝f��^�� ���w��&��p(B��[_��5�4�S~>��F�Lm��A="�e��$j�������OM�`�#�gV�"������s�ߵ2�*k�~9�'���~�D��6�h*$k�*>���	|����mى)H�G��*g'h`vg�2�2)\E�	O)4��5��2��\s��8��g)�����L�^VE0E���ƀ���EdP�e��"�/�� ��s�1HSG�dX$)�� ٰc?&,}.���̮��'�{���+���D��n#�b<�&p�XZn�;UAV��FY��0`��d�7�up��/<���p����8��vh��";�g����R����Ml�f��I��p�R���̏Imd(/��ǻ��euD=���_P �e7�ឺ#���<�q��g�Ggm�3�{v�<�ca��h�y���ks�i�drh4)���!tXcC+��*ҋ93�7$�c�TS���A%��	���������/1�NWi�IraQ�`�.t���7)=��Js��Qa�����-�j�f�"9�-ݴ�բ�r_�v��l0���$bsױ��$]�gz�`P�"7�|���>���x+�qIקB���u�q�l�%;)19�FL�g&��ƍ��>ps�K2M�*�F5�	cf7��ߖ4�D{J�
�k��7�
�_w# 69�X��@��U�4%]���&���t�#o�Cw�1�	x� Ar� ��rl�}0�ȶ#2���A-u���]	-��=�#�ǿvF��;�᤿f��K��UеRǺ�ث��vi����ݼxd��̐�)��c�r�͠���B����:�i�_B�s�Ѱ~��WK�$j'-�����]�(=�@��wL��$�F�%!�$D�4���69P��pI�D����,_���n�1}���?
��O���5�Ckm��wf٢� T=��?ބ�#ް��Զ,�R�1+og�8"�Z�k�+G�J�
_hA�>A+�4}���bٮv9LG�:Wէ6{��l���X�I3�������VM�ק}�e�w�NJ�V`㘬ڹj,�<#e���H���U�*�2\���~/����"��.!��~t���O���Z�i%��ט]�K��gɉؾ� �ӻ�;�L.!O3��͛+>
Z2��7����	M�<6�m��#c n{�����$Vg�(ؓ*��Z��f�
�˹�F̧����o{����}f��OH!R�Гo�X�s+��Y9d�k���u6�R�kp�-i���I����A���+��j����am����@����n�? �e��;��qQJ'�baS��G�cO�5����'���7��sp΅�^�_]�gu�����aX�eA �+���&&O�Y���w�8Jhe�o�����s9�;�a��A�~c��ͤ�L���N���>�ޟ|8)�ʵ������U�=��0dw����s��Ӧ�a�h!�e�-���<0��:�>y9�s�U����F;�|a͸l�9��o^�]A��K��*c,�̤Ś���r��Ai����,��*���r�ٿ�Á>�׌s��9e>�Mm�$�gC�r�`����sV+ɋ�U�{q��V��#��C��2�@�)��I�P'+��պi��-�@='s�^�7�%o,ٔe.�BrC�饝���~>�����&hf9�������p�4J생��>�F�ɏ�Ϯ23V�U\H�Yވ���f$%4k�D����`W���@δ� �8MA�0�Ts��5�tR��Vwa�X,���t�r-�������z�e"��,�e[q�]G#��9����o�z�/@��:��c���!�/ݍo�3�v���=��WSpѪ��W��J��]ż.~�J��A"�7b	�J5�R)��sN-m%�WJZ�L�ͩd�U�yª �}���4�5�龍��D���]��p?G�\�� �E����Z��N����1 ���QزJ��9�N.6���-��0pa�:�G�)��:=<�q�a��.�J�=X�9V	�������*�D�g�8���+���^s0]�[�y֡Dg*�a.t�8`YupN(:Y��^w��@��F��H����Ъ��0�.�ۚ6dq@ R�딇tA>�v>�����0�~�tg[K�-�P��B~�Q���e��t���q��:mT�	mA��6�6�v-��Hkֽт�y�o�{0�p�1�6���VrA6�lX��)⴫��1��uzԹ�+?`W	L���BB�&vJs�i���4�ف�?���j�u�m�c@�2y���Ƞ�`��әL^�k$��Z�O8�$sP�آ���~_@��G7�D̄|�B'�hV��A�a����������ݢ�ô�r<5��9��:N�*=�lGR�$캳~X��T�.�$��4@Y�{*5�!� J\2I��ۈ�;�i��%�p���Kn���r��3��X����a2�Y�+x�{]AC����.R��7a �%8ץ`��S�M��5ϡF@MZw0�K��>%��9y5��s�5\�#�k�T!	���O��ٓfiP\Iˎ[B�������d�ӊ�T�!�9�x�	7]����{�#\,��y���r��l�q�DJ>�n�����n�7��n!^(B��N}��t);8��y&/���"��~��}��6�Mh~i�ܢP?���d�m�Sa��x����5�zO�* �K�e�.Y��&����ټ)"��h���3JB��P��9����Ђ����N[�HȀ���Q���u��:��e��  �v� pq����t�r¾y̱td��,�64v'���k�h��u󡓖�$*��?�+�����o-Ԅ��cO6��t�����
b�W��[�8�J
�QC[��=�Q4c#1��L ���Mɡ~E�[l��91����~�Y��ai���#�(T=���c��!4_�w9�T�B���{U�l�z١:	1P1�9%��s�8�O_���~�HӺ�=@��Z��b�V�A��vW����$j�H�I�I���IW< �8:���O&gA츓
�����1���懆�aq2�Y�4���1���P�*�Rl�`��]��a��H�M�a�i9�gI/)�
[�=c��bD�U5�R^��J�1�!��dH~+�a�__��<(��j�,^2;[�B���0Btr���~Qg��2]��ʳe�����'�[�/�`s�r�a�?����ٺ�4����
��ݘ��\�I	��=���D7�y��2�+�Ԇ ���y"e�X���̇&#bYUK�U5����@�4v��X�� ���B�}��M�z(@ �>)�w#��.pnYB\�ۏ(2��0Ad>Y/�1���f��x� ����(a,z��\��k���o�>���/���خ�q"Lp���n�u��2�o@)����Ì��NTe��a�I�'h���9��O��")���Yt��u}`,,�.)�K͒J:�+:.j?�$�<�&�Q�)�O�#�XSJ��s�-ʓ@s4a�0��K�����p3>ob�`r*���,��l3�.��B���,�D�Y��e�l X��kV5��o~���+�,�~3�џ_
�K�8��G�h�0��aƛ����ڂ����0��@��u���h�>Bx���ՄΣqY�[�P�k��|�!�*g����>�bݑu:�lS��N��[W�౺	�ɟ-�㼹�N<��A�\$��fDǱ[��Uzx.��Ƣ})hp��ܝ��ȟ����ID*H����y���;�5}�{����*:4��M,�t���H���!A\"����lB�-������Ex�O��G�#�6Y.nܽ"O�Zz��(#��~�D	l�,$$�g������L�cm�ֈ5À�����+��@��>(�R9G�c��K9PM�z�b� YǊ2ؤD��YF
Xc!%��2������Ee�=�Y�t�S��mp�ų��!�����g�H��R�B�tI)�Q��U�2�	qǊY� �t��H@'Gܮ{ٶ�x;_��h:�&%T��3�i����Ç���=�`(����7ӌAB������p{��' �����OrJe�>�H[At��PM�by��1̶�D'�"7�R�����������3�J��R��`�-@� _n�j͔���44
1�+&x�hI�2X���A�2[�B;yv��p�Ht8`�V:?0}�0c��C�+&��X4=\Cy��[��,bA5*��nS�y��)����V>A���&A�f��L��y�p�\��*���f���E_���>,M� ��G��gTq���²yO䫸ˮТ�����O�(�)F�`5r���c��l�ds�{Q�A�d����a�)�Y�G�v����u3���f:�����Ug���P���V}k}X�������<�&Uo$���7`5�����Q�fA�x�#5��|V{es~�:����O������Uٲ~�,������/�-e[Δ����(��<d;��(!����R�|k�y������������k�����]�?;p��]��tG�)>�x�Oz�h�p���9�NÄ�1���݄b�80@l�i�"�Ӻ��-e%���7G4���BKxV$CxI/h��,�Vb�K�TR�Ec��ܣ!$R��r8-sv9#0?�,�S�&�>2��P�q�!�y,r�9��$�tlZ7������q?��Ϣ�:���n�;�R�����Z(�Hm�2#�O�
�T���M޼#�p�o�7:�!T��d�Q6:N�瘩�/������h(
�c��I�����ӎ�vo�O���~b�y��˓&�A��Q��>�p���}�\����G�WTH��	qU��x����{E��� �8���N��0�u���\ā�A�9q���%�,uWE
�h��dg�0��0�}8�2�2"���/д<�K�L�y,&���+���͎N{4���
���Gܫ�P+��x�������~�Mߣ߂�mH��r�M�!�y|4�o<��R�UĔz�X��9=��i\Ņ
����T���mS�=��n+�C"1,Ob R��O���	ʹD�	{�G����N�Ѧ��\u ���� ��َON��3ZK(h���)�1i��^�-pX/��\c(�M�����-��pZ� B���أl��Y�#��37I!����;(b����&7H��B����"u�#%ȅF�4>��*�h]ZqoU��^�6�~�0d>�X�,�P��`u�r8(���SŵggE��f�� قU���yA��W�Q��^���p��M7�(��⍙����j�,ؙ5�mҜ��}��T�����X3��f�j�fQX1h޷���-7�"`gvע[y����͆|��Q����ѕ�X�qB�{������ʨ�J��d�nX&�Ӛ�8|�3�zZd��o�-2�S�}�w� �â��Lb8�ϱ�Zǿ��D�v��pÏ$�ʥ�q^8=��r�=��o�=�����I2`�����bk�ْ5��u��59�]Y:Q�i��o��Ux}��a-��J4.��h	-�i��]���2'�~d�T��j)29{�¡˯@P��n�Ȭe��h�^Ҭ*h�W[���޳�����_�t~x0-r^���X˒ĪNR�����l`���.��b���IA��Fο���{��@�pׅ�0�`J��j��c�^7,pj��9�5� �N�yB�����fP�g�C�5F�'K�Y�9ί������e��w(bF�ң�W@�x4Z�;�<��Aa�r�{�T2v���Z�L"!H%	���Qqs������EXw��$��?�ks>s�ɻ���O�]��)����'�"��@u@�ݪ8_K�f��
��l,̵�C�:���>�ܭ˟/ᅲs�!�����	�~�!�QG]���''�	oN�6R���ZR�8�$=�b��Jɻqx )�ߏ�W���T�8"��2CJ�T=�o&�A���j����Rr�1��XW��W8̘yz���@�J�dwPŒ��-c�bt�y4,���rY�W�̥p�'��a�V����w#�7}v󋕫b�e<~���������yRC�o� n�C8�~��Mn���9�=	�>Ӄ��H:�ڪ�AD2�9"C�t��ъ�f����Cc�=���͏~{#���2ƽ�I��ݾFH����E�� �+�TF��-����}^�9B��`�1���%)���T�x��ɍ����$����l�QE~0����~ ���6��#���I���"��].=qb�vH��8^�5�B#�N{�&��l�,n�#i��:��	l[�0u���u+Ч��t����FH^W=u���l���+��l3C�J�7�y�^GߜJ$&k�\o7Û���]��Q+U��%%�6C�emCы�L��?-��#�w0���Gu��}`�q��O
�<��y��@�=�xl"t���-�>������ >��L�X'4)B�_�w�2~��P�����F��ܮ�GI�2zQB���]���u)h�t�{y���&r�V�[E���xu�ay������D�fVK5!T;Y�+�u�p�*�Ė=�ҷ�
�z(��hh�����c�	,(��TXa� �;���/&��7zu�
�b�{_�t�M��B���"��q�_�b���\�3�5)E�ŇM)s�'��b.Ե�Z%�rvq��#n�����nd������~=�[*Z�AF��ް~�[ެ�~���S1��i;H^ܡ�V���:�����1a`��L���Rܐ�,������Yqa��V8~�u� ��Ը��y�jFX�أ+�BZ@2���e�W&����{t���\�>�����|�jΣ�js���B��>���V:uc��1K��l��(yسe+���Z����S�{i1^}������*�'"��gIYY0C�=�q�]=;�Jq��͟�ಈ�֋���O�>�0��ɼK�@q��m��$�ؽ��	�i��V��Y�ي�S�+�^z��x�OIq$;MH(w=���&�t�
���M7����,
�v���"w�Bɜb�0 qC����ZL�;�>գ.��1�E]0�M���<��޽X�� �ӊ"T2��a���Tb/`���5U��*�R���l�^��%	/F6A���O���8H�فv�p������ްϏ��.g��*�6>�F�]ޝ隸d\Rp#1*z�	o��Z����)�:�hJ�Ȓ��
��R���)q���P�y�6����|��� �����IW1����_�����Z�Q�Ѐ>u5�10�}�J�oB�T��O<�&t���7S��ƥ��b��~�>�d�~��wuR}ǫN�r"q�����^"�y3�a�S�]
�����~p`ד�E�����Ey#��9�ft�������?����+e���@���FHq	�ڰ�.w�iw��<�v�aU�Ѳ�2����W����N���M�3��%�	�9�IaN���&�Y������	��XuC��F�@O/,�s�4#Ƙ�r���:���ɶ�_)ט��h���!E����g�F���P�6=.Xo(���]���p
���>���
_ِ�qy�ї��鹯T��d���� A5��r�~��`�Xj�x�g�C#ő8	';�\t8�n�.�?�
��L9��w	�~U*(Q��J'�Y=� O���r�vy����hĨ'^�]
�S�Ć�D��'s3���JS�r���Mi�l���Q���\Tc�X˜x;�ݬQ�8X�%��@vf�!(�n��[����	P�z��{���!��`�H!	Uf���M�������hS��@Li�[�I 9N��s�*h#\��ŌWא��@�@{�L��鶏��?���h�5����Ռ�+��H���s��]ET��M��ń�v4�����pNRX.���1J������{'�	�|sDk��X�������~W�v��[�{�+�N����Y5�Y�#�|����SD �QYiRا�;@�Ҍ�2�e^�����HY@�۟�!í4�4�8%��6a�S����xi> �[�"�q�Y�*nS��"��6;H%q�wKH�ߵPH�kƏ.Q����{�Q�ˡ��S$yj�$� �Q��q����(œY�c����K"s��RZ����y�Ύ�"�-��Tѭé��-�$(��-*�X�+D��W��P�x2o��p� �8�S�,k!m�����,�x����v�up�x�7����뻟K'|�� ��3���:!�	�����G���;}�#c�*��
>��*�8��U��������a�}�i�r /F������$�uB4j�le�,r���BXX� �)F&�6��FK��ڼߘ=&���8H>�:_1�<�#ݜۊ��L��c��S,��́ݎ�&~��U���_-��ͥ|9^B����ٲ�#��q65 u	/�k2j3�SpS�ێ	��o�:�kI�D���g���c�]�RMr[io��zP'B1�Bj�(u�{�'h��Xt(Z�ef�p1l������j��h�h�7{�h����V�A���'�D�&�k͔ϼ��%��>�	��?do����8����*��D��'�o c����	��y|M��p�Q��N���q�Z[�$9��7*�*�L	����P����Z��=��R����?2Ln�B�S��`�mE�R��`�S�n���OI?{�����>�F���*�+k�w8bGRG��Q��E�lġ�6k�A�)l�/*�3�Y�{Q�qZ;�w_��$q�P�<@�t��P���Y��zI��~d~��]ψ\��
4�cW̡�[��6��9eOb4+[��ʚ�&��Z� ����*���3XʢY7><o�4#��AO�!�㻦
q� ��x��!��|��<��I67z�ה ���l�J�Mꛈ
�jy'�FƔ����c]�e��\��Q�Ā�z���ꔬ(�&�i$�v���?X�s��ʸ���7�I�W�����pvs�~��_�����>�+ʨ��>H��R�.�nĝ[��o&�7���#���Q�c�W�TU1Q��B3 Q�.@Ȓ��H�Qu�Jʣ��d������ek �ω��u|�f/���:�������p�1��q!AU~Hh����$S���Uc�'�9Ŗ4��tg��ϳ���0쭅�*�����*��5�R�Rf�����Hִ�Y3?��V�Zh�44m�C�	E�)�U'e y�o]�\�Yԡ�~7 <F_)т�=w�Ӡ�5����H�L�K!��?]�ڃ��o�M�DʝtO���u��m\!XqC7k2�X� ���"5e�7p�d�c`T�)���3���{�(<��wS�f<L�(K�] ����N�*�ĸZ�s��A����{��jo����%,��5�{�	�̪������p6��x�F�<����/9����U�g�D�}ؠ2����n�y�_c�y��{M��[1&�W���Lw�ZM�d��oVt��F]Q����%{�%Gy?u�۟����b{��cu�v�3u�	�����<M����@�qZG�Z<�Z������,l���l��-aE�`Ճ��F�Џgâ��Ɂ�`1�߃Բo<���.i9^9Xt�1��[�����@�'�6Ke�̊����> ��S�q����z�����p�پF��T[=��ﮧX����2���H"���Z@]���'ܿ���z���~3�(�F�����[�v6�A��z亿���׳�6�C�.�M����Q����z�}���P��i��߷�L��3Rk{Or��{�����QC���է�ķ��*�21q��`&#�T�ҡ�53P�^�q+���9r.��T��)��L,�h])m��Gh�`����� '�% )��T�'�6D\���t�+��g4��d��G9]ph�WY
<c�v�?��Hg��"���td��oF�E/��|��2S~K�Tޠ��H��$BY=f˘_�h{}8��1�\	<�� �<����y8�{�dY��p4��6>d+�ƴ��L������S��:k�=?C��.�^�)��t�ȴ����	5z�!�4YQ�!�;�a�'�h�+�fd]C�R�ʏ���fLVu�$ ��BG�1�s���?�x4�+�GC0�^�/,(�����$H %R�\e9mf��ٌ��R}�m orJ��A+p�6�xk1q���*kyB�kVE��"��;��xe�l�Z�6
;Ԕ ��ʬ��"��
�"�1k��{��(*F{�����	�{q���e�Tz� i���
A�q��k�6�%-%"��H�=����Y������Mg�Ń�	sŇ(�t@�������jsIM��]̂�7T���:v�jCCh�58��@�� �E�.�	NѤ�OP���*��GV=����Cv�]��Tl�*�˺��N'[��B,���Vt}}��U�3-΢z���6���/�xU�L�M����/h&j�,^����*E<� M�+�[�Y�e�EzoM���9�\��J66�����,>>dK�_Ȓ.��o��rLO$���z��'@Z���m oȋX���7k[z(qP��C�oݪ��pP�W�]gS�EB0�!�� vOJ�����Ua���v_�?s��ړڭڔ����Hf���o�w�b��QX��\i��AD 0r:`&-�����aMr^����`��:R�6��%2�� O�Ovæ���O@��0Y����R![�.�ǈÊ��,r��+�6��6�s%�3��VIK��E>�v��H8��x���Q��-�e��0�7�#��Ø9�R�� zwX���b�Vk����9�7֬V�����F;��ҽA� Kխ`�~;h.sxD�N	M�e�M@����#^��79��$���PWܡ ��G��W�DMz���� ?A�"����м3o�����Ҙv<�l*�0'��G��В�C胧�h#I|�rͼ��aۢ\erR$V��i-�Pi,�[i6_M5�![׍^a+=�=���剻�H�Bx�^��Hp���gu#�u�9QZ��h�)M#�K�VO�K�/RV*]�Z��s�J���bU��\��[�ɛ^��\]ˆ�L��F��ʹ����^�@'�u'�/z�rK]lO<��.�+��^�Iy��� ��Oq�rSD��8T�)%�S'g
W���/��E�~M��HI����;�"�X��qŴ�fѺ%�rfNk�Ƈ�#�Q�*���ͮ�Ş~l��Ѓ�"�@��@��2Q�+otZ��@nKผ;�m�h�;��@�>��OJ�m�*6����> ��Iw��V�36�ϱ�NY��N�ݮ\��R��&m�vK�3at��W~tt�z�M�{
l0|(/5����t���=�ڗm|Eyͅ^�A��ulk��P���Y���@/51H�ix~��/�=�m{g��"�7 �!� �a�,GS��Ϣ�����wV�A��0ćZBh�t�ya�\��X�T�7˭W�
P�Q�PYŷs�k�x4�u�j�D��]��~�g3���ZG��Y�3ao�g2#��KE&b��ŭǞ��dMV�ˎ�����#�!Y_��M�>�: �/,���܉�\���������E�G� �֖���1J^���0	�[G��ul����	��	z��ľf�aڹ�JĐÌ,00MY8A�k�(��b�����@Uw�^����ɈbS�A>�ƛ��Ǚ32�k|��Eo��.�%fM�|��T8Uc�0Z��Ŗ �ț�Qݛ	A�OyL���^�4V�Wq�[T��.�L���]z��Q�����p��L ������i
jS����IK���0ʀ�
��4�▟�
aŐ�dŴ�,4�b��Ȱ�:BA\7m�����?�F7�u�E����)�
~x飙eE�OJbr��|U��k�&V��E1�o:R;��Ȗ�:^B�4�F��b�ʠM�1��ϫ������W}d^��(�K�4��_E��݇=L/�ӂ{������Ec��S2�����"��$q���Du��F��/���~L��c�e�����K�C�@9�.ˬ$3x�y$(&��3Qӽ��V���1���G�4%F��w� r<�/�DW���7��C6G����U�_�9hcxP�{;5ꣁh�A��cT�ޮ��.�Ѱ���g?�({�F��Qۼ�Zr�E34�.�����T��JJg`'RdW��W��͏kZ� Q����ɱ33�~��[�L�]����r�����u�_���X�.ͼ�|�K����ۼB��E��m���R�.ȋ<�&�3-�I3y�9cxh�d��4'u7«2����7�;�#�y���`2��Xdx(q>�h��R(F h?�6	�)fҳX�WDZzyn��=���G���2>�M��0��ohG�V=L����g�w�c}jL?�#�*�Q��iv���e^X�R^
�)�%7˸�����ZjF�y?�h��y��*��
сjc���)���Z�TF�z̮H\#�s{ϟ<1r���"T�;βd?(�*�\{d�R�B�A��sM(�o'����eMxY{�JD�%U	���0��������=����<��C�K��sx�p���g�fה'�KX��u������(!𓢺^~`�n1Ǚ*�����~�u��l�t�|b����[��;�ć��*�k�\��پS����nn�.�fIk'D��)%֓����$�j��u�s�1�&�r�ZM&�j�Y[�k���0�!���h�>���$�#��W o.$�hV��zNRo��{��a�;�HL �@:F�BQ�vr��?�<�x�(
)+�"���!������"q^j�v�粔>(�PC�����D��m����K�Q�.�/�UTظ�a��"��7|�Ȁ��!���aOg{�oS��*�'�ӧsU�l� 5]���lb�:�Pf�mG7,�Ug.~=��8�]�Gް�� �	x0�)bIO�5�:(��bɊjo�E����1���'���5/j�F聜���HY�����?$��r�\��?r��;��i��9���Re��D]�Lʀx�~l�_@뺫E��� �I�)�(X�a?'۷��s�ƾ�(���Y
����駈xD�f R;/�M<�=H������M�CcȀ�L��(��h�i��Z��3-�ܒ��{�s�����6<�O+������۲�9������-���	$[s[�>�	�e��¦&IM���4ZT%�t�������Z-^}���G�����:��F����$cHC�W�#p=�>w�%u �� u�@x��Y�@�k3�)��[��I7�A4��:�X���x���?���{"�c��7)l\�CJ���_�C�����oj^�؛�#��Q�S��m�J�sQ�`~K�k�SPjXqx�O�f�Xb�C��H%�x
ݔ[���n��\�e�_3c4��2�"�
1o�ׅ
�ki�s����(>��)����o��6����R�F��<EG;���~�re<�y,�}Y�n�=�4=SWa?O�0Ht�J���]EG�Q�hz��|�͗g�����je�F�RDӢ3^�{��Y�Q(I���.��=FoL</���#�	v���<2�)%��?��r;�I��)r��yANIw���@�?͍���kv+2i�Uk4��6�~s�B4Gv�[�� �Fu�!k�����4/2f�,�>��wܹ�-�)��服̷ p6
��'-ɩ	�P�[��^��d_2�3-��d���`��a��W,(1����/���t�x��T�K�G����#S���,3��r�sT}آ�yi�Y�(gw�k���#+��u��,1�1Od����<�������-˂"��WRcLBN�����5ж\n��G��0�B'D�Z,�g=\�"�g3֐arӞnpSP@m;��V�X�s�m J�-��xkw����6΢�`[�u˞��^^
��d��pZ
&�^����}~I�&9*��6sΎ�|PƜ�k��A�����Gz!5U\E60*��
x�w5x� _2�,zm`+r�:����ԁҺ�E޺m�j3ʰ�ߪ�?2Ӊ��4��Œ�>i�ϯ�Ύ���#�xa5�Y؜����kf�;�r�Z)5�N���,xD�0�����*u��7��3���b=�y�N�k�#���%�x����-2�㎱tm�ǫ��(Ԝ��{�����ߠz��+�a��}1s�R���?ڻ�g��a}աFm�����HGR|����檩�G��p���sh�UGXQ���,��ƾs�y^r�I�]7bPL� RD%A6�Sw�E|4�n����{Pt>����^�Ԭ�rɝ��f�"���(%��Kd�W��uɺ�߶�#C��#�P����S�<u	�&�W����D��nM~�X��:��q����t����wH��=Z�Q����f��y'iX5�Tozvۥ�h����B�:�e�,GT�5���D�i,�%�]�m����ַ�[V$ˀ�4V�ʻ,s�=�|�_��3qE�$��A'���O��kn����PXJƏ�v�)��z+�$��d�w�:3�������º�}�tc�A�����g}0�BC�ց�j��v�ܷ])��6U:|PN��Ӓ�!@B��9�}%h2Mx����ٻ��84��eT>�p�*A�P�;�����a"[��h~��D�����VN�Oy����E��������$F�9��� &}��
����sS3W?����.��	_��yOd��5)��IB��x55����׮{�����H}B����˰��̙ds�@����ށfv�I75t6�o��-r��˜������}�"yy+�]U%�^{�Ӆ���ݬ_��I�_�6tWV�M��Zv��eh��Y� E�B�D���'��E��a/� +�9�w5����26�ҙ:p����N\��;�VP�y����b��֚������9���u��j&
F�j/��#e�f/0'���	���I��VTO� �\�Rܽ��<		c�'H���9��L��"��!���K�N�����b�X��'"��U2�r��,����G��,�O�I���:f��r�r�޺��<������`'����]�5-��Ùf���ⱘ~\p[E2�G����{у�Q��p%�Pq��5z�m�=��5U�=L��Bz����zx���1t�l�"�Qh�HIw��*|��6uv#y���\�5���r�v�`�t�N�����؍��l���)�����,�nB�?�8r<��@8^�?����]���~U��Pl9 w��G����i���UQظC�' A-~�a��X޹C��}���`�S�Q>RJ�h8�F[NA��R-�rW����-6�|8_��v:5@]�#V�`H�
^�Q6�8�y0)�=�E�{�ٸ$;��p���p�G�]aG�ܴx`ؿ�L$b>�>)(xȾ	99�3�M�!}�r�uN�6e4��}�x,ٚg��;f�[�.N���I/q���V.7�[��Gv��q��`T���}2%E`!�!���U�,s啠�`e);�~O`�wT���PHp���\���M(�����X���s�ފ��PU�����_D�w]��)q�T�;��W7��f˪$���X� #���a�K<�Y[��)�����7��a9� P	�*�yBTT I[��p��y�OG��ў����A����b�������2J�V1k:�-S�
x
�8>�)�˅��+�!��j�ո�"K�=��B�
0��;�j��Ӧ�v� �g H�n�N>���$�9>׽	���jy4H��ϴ�Z �!O;1/������0�>ǂ��3�6b	V���\.M��,�p���=����bz ۛ��>���?����3�t���O� �i�/�ʳ'JWpt ��)��o&a�Ƒ��.X�ϐ'7p�f1R�:h*�hk�)���������g��-ʝ�BT5!`�h+x��g���W�l�T�ɳ����6�5��>�k^�y�;��Dt��]����VS�e����f���/���pEN�����[��4��鎪T��hl>�Va>6����BW�`Rm �K���� �Q�p�
��n=���$M�{�l!�̤*�gboO:����Y0-�?}�T�!��\w$�̥˵���?�<�~�[���8���Zf<��?�D�v���c�*o��5��"g"el��b����~s�g�#��ߵ�o��P9��<�z�ό��pz��J�� �p��Uz�M����@ߏ���P���c(_sn���=?�4�{��ax��X��4��AS&���ҥ|��N �ڧ�^�nM�'\@�&/�'l��'`ip*�F����fġ�X����jgodK[���;e����B�k�����V�-)@!�Z�L��{�W��\� ��W7 �LJ?y�QI�;'�<�cj���LR 'Ɣ�����LL$Eyѳ�*z��tf3r�
�����)~�]
��(�����6�j �M������2�\�����0ӁսZa2w��$ ������'�����n����u��+�ĠD�E"Ȅ�~pZ�P�d�qy��Ȩ�:��ΟXе��}�r�-�Оm��Ϣm��s�&g�&��cv��"m�Z�+8�^p�Gl���� ���|ʰ��uK[&G��C��>���`h�%�e����m�o�d������Z��d�n\�衦����o ���&�w�,�6F&�!.�=Q7�4v���w�e���F���u!Ѐ�bw�ZWMgdG¢.M����uV����	͆����N��YᇽX�_
�6���ΟR��~R�n�a���i����~�H��mb �p�]I4z�:��g�k����A+=b��&(l6y���oxc����+"�'�i�b��RҔ^����Y��粻iA���!lg��0��z�MZ��tk���
��E�1�<U@t Q�vO
w�{kL*Y����^�oyuh�^㉤Y1K��m�>=d� ��8- �}:����;�T������q������AکL�d�7>��#gw���\�K���y�#��h�<딘>]�C��B]m�>в�O��ys;���#�3:�z��Qs�Q���]��7�a�����	�6J��0�4]�ϲs���2/��[>䕜X��ׄ�Jm0gp�ћO
�����e�rX����� _�J��ѳE�0�t� �7�ܨ%�ፑ�XO@���H�S�m���W�Q�ۣos0��e��'�`���G3�����WGBa٪3"��������Hǒ���4��eT�4� �=�j�I�^:��ŭL?8���aeb�.���X�I��f]h��2rr���\jqR�<�B��5��&�|�ַ"�;<�-:�\��9�]��Ic��kF�<BT��j�!� jVIvǛ��[V����oS�~�3Nw�b�ܬ���� ���d/���=����I#@�
���(�~�n�z�A�K" ����c���kpx�ew[�N���G�6i�]�:�0���u�w-�[���OA8�/�'[g��Y36iKP��r��ʑ��'S��f��t��:��#�cd��2��&�_`H�	�b��B�x(��<p5L2�}�摽��k�a���8� �����ԬEh
�a*�#��B��/ ��/�]���>|QT�&�����/�����(��Q\��Q�&!۳�����Bn/�R��lS?L(�t��:�������U�Ca��\n~8�
�ƠP�2�:��-��@KN�����h��n��~g�����x�u�Sw'O1\��"�{����a���{Vn)kK��`IK��d��n��̨�&{-z��rK9��@�W���I�ۖ�4{�~T�n�~8����|��x.q4�e�MDIÄ�ui��E�۬�������xQ
z�G-�}��8BA%z�Fr�n���#���'��9�1�6�F�|M�B�����-o�{���V� �����o]zJ�i+�|�{:�ɩK�����5ƞ:�#�q��c��8�=�B��ad8ܱkbJ����y |S�8�����6Ċ;Q*5�N+ᣳ�#�>�����]�4ꞂkHع;������Q!��fĪ�>�v�Ψ��Df\��j�`��k`ğ��'��VM�����Z��ڀ���Э��|ӨJʕ��_��\JLxx(��iJ�&lZ9�k�2�̄�*�툜�f����MI0M0�}H�.e_�����I�E�n���O��D���Cv���Pl�=��Fk�u�IN�b�kMY�WԾ\en���i�v+�9�e�_	��PFS22oT�x'�����t�b���C,\�9�`C˾�2�{������3�#��;I�����p���I����J�d��t
k��75~X��]�0u��	��_+��k�� ���)K��wͨVA��'���X��w�����@o�SO�^���Nb��P�Y�xι�*��T'����#�S6�{m�N�t��F��=�aCKojܘ�x��"m3?�0�j����p�0�V`7�e�h}*4-�>,�OSDKRYGWKz"N�Z���"�p�^�^zn&�A��h�,?T�A��#b%����B��	���!7Oh!|Lkᡰ�ҵ�=r��Ke%��v)nZG��������CP|����wWI����
��SC��<!���+c��@�*W߷�=�|ڙ�LX��Wxh}�B4��Y�뚣�@9�[0���`�ׯ9[L����(q�\�~Vм h�TM�KǤ�1�s챙c��`rٔ�.@|������ʙz{�&� ��B�x��錾[����k������hSՃ�N�2h���;�!� -fȀ�a��^E8N;S�Pt]|�0�)L�˩V��q"�FƔ��ɘt�ҽZc*"�@��~���YrOA.Q9��@�Ë��H��W+<{p�uI�ϩ%I��ʁ��Y��؃n���M�\Sɼ�+�Y�\�]���jre�s���G,#��-����A��� ���̥ɗu��oJ�`j��KvL�	��nS��
A>o�2ܠ�]��"�*�6���ٱ�a�no�M�˥�[+�^�1�H���5���Z­��Jx�L�Z����!�6-}H��BG�z�W���ރ������'{j1�y��`��V�f�e�P�����^Z�"�[�b�l��J|���I�!��%���L[���8͑:��깈��UP�_�d����?�}:90{2C��$�A�k��w��L�9zMK1�
#�V!�:�Ȉi�2r��./�z�%@H��
d(�ha�AR���	b�保@��Ղ��������.� N�[ĉ��o�|�Q�uȗ.����>=���-`�F挫�_
��T���X��$^��S)��b�������������u2�#���)�>r�G��CD,���P��!��ʻn���	:�@�\�T��x�������������ĉ�~�si%5��"�LU �;";�9P�:M(C��,��o�ǈP�ﶹW�	ˊlQ"-�k�w�����9܌b��/���;�E/P�EG���U ���l�v0�gL\#����nk�t��o`�v�^vw��w�\ L��L�/V���w�!��U�w�"P�0��ԩKĀ�$�ؔ͑?�'ְ�/�^��a��$N��zE���6�����Z����Ɉ��uw_�D)����p�!����J�fs���K~�K�^w�X���:�o���gK�!� ��ك�Z�!��Q�����;+�ᴆ��u��MGy�:<[fFaݯe�"ɚ!j����Y9]��������L�f���:���+G��s^���&|ʤ�u�����+ �(
� �пP��C�j��ݠ�:�A����G�T�k=�������^G�3\Z�"��R�i��H�D�U���������b���٩���9yVr̷���ߕ���5�r3�0�ʎ��rqٵ\IAx.��"QR�k��=��"M7��qlxɿC4o�^����o����>�Y�Q�
d�ER��}���x-�},��o����q�^�%�U�-��\�3�X�{J���ebP6*�ٚ�<a��jy�	���c�uĿ��8l]�Vi�ؙ�]1��B�Kq�Ľ�Yu�O���B!$�0K���d��:ٻ�� ��������Ec��kfR�hU�Z�3��~�n52�v{xGzQ���%-	��Y���)Z�t�f���So����f&�RQ������AW� x_���4/d�>�11}4ʹe��-I=��-l?]���)ph���&K�qFPN��(-�M�r
K�$��>"�a�T��T�ᙥs�*�8�~�G��h�<5���owZ
�wz�h�`��
����r��#�#X_f�AwTs�����Uj@Z1��h�v������[�\�y�D,���Yg�)����|�<Z� Λ���03�.���eG%��$>����*-��k��x�"�[}���Qf\,�{ǝ|�QˑaT�e*{��7��mDR��l�QH���{T�>���[�t�F�5�6���M�pAG>������x����OQN���-#j+�i˹�ؙC)��q(� |���1�i]��	j����F^��g���f�*dP��̽(�έD�\)/b�b����X��߸G��g͘�E.�_�v����w�(v�,�j-��X�̜#�r�Cq��w�z.	�
:���w*�S�~_˶[&J~������JR���'�V��P�����J���NȫG��Z���+F j騸��>R�I�������pI���n�������9�V
���<+���"��)�y4�<�\q쏮%+#�z����L���
9���"Gh(�9������$qYp4���r1�Q2u�	~m�r���8h"Q\��
(�[�ݳ��e����]�z��ծ�[�S5H�����?%ı:m��E�b���9��Oa�Xf��Ă;G�@����A��ݭ;�4b|[��?���B���y	Y(I��{-�TWG���x���+7V�8^��](�a��G���;�G��@O���n��/'�9�:��$�>0`��R����e#������)�؈�g"����DU:�_;ݘ��*7��ƣ����e|5a�ޘ��m�$�+Ǣ�E��y	z�b%�����t��E�Oa<M���dR�59�Ck��`$��P��YeM�)Lm.d��T�i3&jD[ ��@ȍۃV�sWP\Y��hD!�r/�u}�5,|)�̟��O%¹�lt�,����"r.�r�hɺ�;�'9��^&��r�/M�Ji����l"������X�Rad���m�"
)�� �O-�0�����v
�R���U�?��Y�(�=4Bs�.��:�ۊ ӢO/��%�F�֐�Z0�+\j���	�;��'0�V�� �^�*Lo��}��p�u����|a�d����8���RJD��l�h�$�h�C%����̺.	j��??�~=B��xj߃m}���[�P���4�9������O�`
��|�[vvae�UVR��k�w7Wh�~"�B�V$<s\H>��b�;?
/O!B}GT�a��e����[��T'�>$9�k��|�+˔��;%t*�0����p����N������l��y X���꪿D��n���������}ñ�d�|�Д�G��Q��J�C�ՠHG��]�C�OH��hQ�I%Ԣ+�sGm^��:j�^O���ʦ_<>�[}�t�����v6.א��w|D�I��M���Y�)H	���b�}�c=.u�<���o��S��`��?,FYc�,��c��u���!�ݏ��[Ҷ���?�v7S�?*$Í/N,���1��%< 0�����yȡk3n���m3�Wv7�/�^1i�T9o�Ts��!��6�:�{����J�=��
���廋�w����t����m�T�~����5S>JuMva!MG�,����4k�(sg�y������F�"�d�t����N����.yA��L��iE^�6j9�'�h$��*����՞k��~���X�f�m�\5(�J��՟��
εD�����w�dT��(��[8]�vYn��=I����\7�F	O��A��3�eUzz���P��SMB�oXUŬ�OۖC���p�<��[�u%�v�a�q����tf$��??Y<J1���zy]�⡯Z�P)���<gq^9܌WV�����pO��!o<�Z�Ja��X�桲l�a�:�	p��q�0l	�^J�@��vr����=�E�Z)���4 B�Ċh�inVV_�i��ڕU�G�q��#���d�ki�W��Y2�'�Ya7&gE������'�0�
DXZ�i����p�񙕣Ep
�=�:��l�l��h���ܴ�fʗ>0����ډ��=~},��FWl%��`���Μ`�hOY�3�X��Ք�5���[@�b�g���ݣ�D�/�����p�
R�O�/���j?���R�(�6e�P������m��^}���b�Ӊ;�"F2u�����}f�v$Vk��Fx�H��K��3Xs
�f����������^1���tJ^%�%ˡ	Y�z�A����d�����I��,C�Wk�	k��L���߿�0���.n�"S�/A,X�����`ń��#*��3��a{']���7+rK��y!F���!5#����j�Gzb�G�T�G���RI��@ݣwt�/ba�"�?y˽�>�Y�s���f���Ap���B	��y�)9'�-T<��#�n���Lt��B��b,fL�Su�0��)!�O�x�]K7�ϲݯK
�҈�8?<~�/Z*�J�hPӹ��>l�"�巯LE��d�VsÜ�b��S
��j�p����>��[ҵ�_D�P�j��Б *0\>2��Ni��ǽ��و��H�L~!E��M��"������VY���.�rQ*Aaq�NO��)_�F"m�~��,y㼉�� �U�����'����$�@QI't���t����{�X9�Ϳ��А�cv!���ȝ����V7��՘}���G*�������W�O�ܯ�l�2�ke�V�Yt��
E[��Ug�w-��S;�y@v�7�w��񭖈�ӑZ(�-oQ)�����ݏ�Vm�5߁���0��:�d �w�bDw �`�ɴ�LS�X�8�o�?Z*��R5PH����m=��e%�>���/RTD�,Z8��\���_�^+�i�*�8U"�Ձn���/��j�D'(G��$aƤ�p�N���j�;�ɐc�-�(B�ۗaM<T�V"���;ʞ �l��ؙX�̷�L�v����Sy�kH���!W��q�=hz�p��QQP���Wx#}{�����<ޛ��r�u����H���u�,���?�'9�3,5_���S��1�)HD[�]-~����(��$���|�ف�p��v9=�< �q���1���-�=���v���6�|���ykO�a.���;�sPp��z�Y~̿����[wVJA��bg⭒�leYl����dw���0��7e��#WE��HG��X��Z�d���u٤� aFr��4?ظ(�{�lgã�`����+��/=7�Ȣ*W�±���z$9�C��~����b�y��^�OE��m����B�ˤ�+����р)��k���	lo|�0�M�+�U�2��4��#�1�ݳ�e��M�,�Z��t #ٔ��wф�ظ1x� ���t.IH[Kі�VG`�KG�t��u�R�<)�Ü���_0
�Til5r��r�(iu ~����إ���}����? �6s�wf�WAUd#�f(����3�����dAٿ�h��:�jQgӔ��x ��~�9��,�J��\~�t˗��I4f�{�N��"�ⶫ���N�/���+<����\k�ǡF���(���^3�����#��CCkI�3{��������e6Rз���2k��]�j�P
E<W%|s�9[PBe]<{�v��?U<ԛ�NnX$�m2������Ǳ��a�^��lr"`
�[�T�9��ϵڡ������$���"l�(��?��w�[<���]���9&����2�=�����.�;���F�{�Z{�(m$X�L����F��q����z����!��zY ��[*�Mc��8�cC�ٮp���Z���s V+-��oʽ��_͞��1�G�MD	�W5����cyt�]ݠ�x�TK9�u����_��vo=�$��C�a�k�x�牖����F�� ;�[kB�yA��O��������/Z�l=��Y�e�#��4ed%Ŵ�J��6LZ]�8uP����nb�T��(� ���p٢N�0<�f�֙���S�����자�x��~��8l)_�{ܻY�%n�o �[�u��
+���h&!'
kGn;�\����I�qs����Њ��$٣���'����`k�D��JcC);�K|�����Rv\SJk��V��Xe�hv�d �f�R�7#سY���>Ai� [Hz�ň�;���a�*�"�,@�j��Y�7�A�J:pҚ�c�\f<�&�	�B�E�L�R�GrP����S�N(΃^�}W9]gFQ������[��;���!���`����Ʋ*R����{[p\���{�b4��mY��c�$�O�̱R4O�G���v��p�5o���:�vW��uGnQ����N�h�%����s�٪�U)�q �&�7F�5�&"]�㫙\9��j��3 ��)a��\�6�2��� �e�`4*�ysª;@^�b�=����R�Ɵ�L5�}N�>|�ߚ����¤�vg��[���k+���{�.��prc�	:�A�@�E�|���%�8�tp����E�������t(�x�/��5y�"�(u��Ϫ�U��Fm�������)�������Q�$�� r�r�/���Q��6�Z�d�A�%t����}����vʚ��8����DgFg��ce�v��>ϡ���P�T�m���l}��������� :���m�ƞW���!W����W��d	);�n�
W�/����|��U�S$�-k�,�4��X�F��Ve�'ط����v��R%��[�k�?J|Ԩ�d��-c���:����B�\ty�����:Rv��T��(�V+�i����4bz���[�)�*�%D�o����Ő>F6�혜T� hJ���4��XM��n�w~���ћ+]j��d���S��Qc����$?������$B��Y�P~���|4@5.�n��u��XY����T���6�i���I?7s���9���ڣn�gu��:MN(`d�U&�{��C�c�xc�B�N1�K���� LWrL��25eSE�q7��Rm����/��nF�Dt[�eH(��h��/��M��	E�V��-A�������U"q��`@u�^��^J
�Ȫ�<5�l�;B9���sYZ!��d]}�����/Y�{E�Da�7�x}����1V�O8Ut�
T����4_���F�>�w��}d']ֹ��u�'z�:�s~�e��3n�)��۳X�I���Uw_���z���dZ��L���+5�/���8��k��\�/��.�"ʸ�[��l���@M�2����ly ��;�g{s�#�po�Lr�����;��������p��zJ��J�󕞂�^����tYGk6��Kt^��;JE��BSf�s�wzC���g��w�Ͻ�
T�F\Ь��l`��	��Whg��������)�BL��W�T$�e[���+t^a��)���Q�{�\���zZ<(�W���=���h�=��A�p+��{�h!y3h��zđ+�E��k]���L�4E6��˲`<t߉�j%a�ŉ��=3 ב���DM*���
n+]�)���b�So�G����ݳXW�biM��U��1����a�����D|M��nw�GPIef|pQ�2p�UsI�r����}������B҂��-���Zr�q9��6c����4*x��!籾��E7�9��G��p����d] ��\H�9G�ؓ8~���~���v�!��Q��p�R�I5���:��r7oļ�S�A��Asj�E`S�0:B8�����ď�A�L�]�-08QcA�B�亱�i2���'�R&?@��	���B��u���C�K���d����Y�8�+������ޘMK�@ӡ��r8�/��؎xL���t��c�@�dc�����E�6�৩�X n_�m������2�q���Xa$�_� `N�y(�i��,ymj�~�$����~���_1��1�.���V�c�S~E����ӗ�|�,x���P�����3�E;�;�q��.4QaoN_�s���G}��Pl��ة�!z�.r����̞�!�~wC�T�GT+M��}���TxV �2~Vʜ��$J_���N}�`�,Wf�8���-/_������a��ʣ�M{E��j�a,6�-
�[jI�N"zV�@}_�
��0��Ah0T�, �0�H���dg!}�ң��	���_h�q�ښ����X1|���ZT����L�;	�������rp:v�KX?��9d#)��{e\��mc���p����-��]n���;�8ê=�M��fY��7ߠ�Nep�AH=��|(O����Y�Y@~��d���A/Ь�FH]bE�7��%�/cY6����w?z9|Z��p�����7�#����4��:_��zO�mǸ� �^��S&��y@\��%�}�n/_�#f��e7W��@#o>�6�G��@�ț��^vb�-��r���g�/���17#o:p�)rJ��Ǵ!̀lsѮ}?�xA
�e\KfZ�Pn)	osQ+��,�S!�S����.�n���kJ����Wj>}�xc���1��6O���o��ā��$m��M^1;��V*����L{r%��x#O`���N>��W�hD��
Bx1U.�(��G�]�i�:����C��D�<r������Ya�q��}��.�����=�������z�#}��Y|*|#�����c�|c����>�v�OB��T�-H�!S��� ����*7�=)KX��-�b�����;��s�?��/�}�alC����&���i�zG��������·y���Ii�S~rW�hm�E	�d���j��� ��D��IV��������j�~C(�^G����G�#̔Y#�Ȝ����T��Kl>G��'��R�qE��ͽ�!9�{��`A�F?��݀���:&��g���H�5�Q(
k�2�La���O �a��ѳ�������bQo� �]��o0c�|mu�x�v�������f��&LfQ�W\��K���g�R,6�a	f�;��J�E2��<��e��"���g��å;])Np�2��S��H% �!+�0_X� ���(�&(��*V`cՉ�b ��	mϟi�@QE�U��o鶠o�b��}L1YvWSq謿;�W��R��U"15��-ͱ�]���}���o`N���ɼ�� oi�T!}v�{Z\eB��Cb�{��p�KW�dଶ���zG�q�Q,/�6A⻉����Yz ��Mhᘪ�������Z^��ɺ0o���",�&�Sb�U�)�C�a��ڂ�H-[��/���/7�����G���3��D�.���5f�l�R��!b����:n{'B&�r����ʴjC��4�v�1�b�Y|X��=T]s�?	S�Y�����~-G"���[iŶ�wԫ'���J���0Ѧ��+��^�v�?o3	헇�ߩ���c�b(�G�Zڽ��N1$p0
�q;�P�#s���L Xh:'`<�z�i2*��}i4w�'�e�Zj�d�rb��+���A/��$����xj`"�������GmM̰X_�~Ք�+�H�\���{����ߧ���Sd�P�$ݕ��R��u��fq'��ᆎ��-\�}n�u �AU�?�[���wm��~XC�>�0��9*��^C>��Bp������BJ{%p��&�ĵ�qZ>a�^�ިg�Z|> !�����R`���#��e:�Α%�TnA�@�m���elfV=`+���؜3�+[�<苶90W��)�E���P���W_v��}ɬ��tq�: ��"��ъ���/}���B��NX!q���s�Ydyn�K[�v�	��#���
e�w+��Vv�3���ʂjb�k�
�mS�%��[� F�z]��rr#3t��eد����P>X�����n���͛U	0N�W�o��~��{`<Ȝ�u�
h 4�������\���_�4O�O�3l5��Ӻ,9�]���Wkѥe��ZT�[� ���8�������(��D�{������5�XqC���ëU�M8@	H�q��l@,]�y����=��Ѩ�&�#�#`��"up�˸z웺��m-�'n�<=9J��!8�y���2@�������==�9�;�SH�pt(rT���Ѵ͢D�2,:�Rp<b\�?��)J��͑,�ZZ:dw�����1*.��S�#�d���m�x�sQ=}�[�Z`\�"k��F |�s���_�aX/������<ƟD��S,�c��t/��V������Ki;�s����,�����%��r�k~�o�)(;�e��Mi�d�>xl1���Tq�G"%���Iyx"=�Ia�g�z��̢ե�IQi�n�Ѿ �ɥ����>��{�I軓
� y��q)P��V�uϥ7�j���m&��zj.���B�@ɔ�Ex���Ȏ��`hQ�xgyAG�\="#2rp��F�c�	HH��8����5���I����j�'����q@D_� �0��)/�w7ʆق홹�q�����'�)�ث�7��0�D��$�4�$Y�I?��R�2Ŷ�jbƏ4ցT�Gi�����A'ڨ�`��@����B��f.��|W}0nٙ9���ƍ�d ��j��T�EJw9p��֯�� ����:��%�c��貿jg4�䉑 {����tD�~7QC��^`LkugK��'�=�eZ$䵻�,d�֢6��j��]����	o�oP	E�.��P��m|�^ a�7t�H�Ę�/==����i���g���u7*]����p+V��U�4��$;�_�ܧhL�}QH5���
L��qj�'7�=��ʠ��VK�����ߓ�A1CRwl�y��jO,�f��2�1�ї�Ry#�����w�N�[����N�?}eL�(���:�@�|�₦,i�~ʳ�R8��N����j{�$]�"m�����H�V��ؔ{�ȗh%�����$1����`xXa��_htB�5e�un8b�Ek?�'n]!B�JN�f�9�Cp]f�H+ho�,�7�s�WBun�����z�^bx��F��� ^����g�y���^,�����܆���ϔrZ�����nƇk����Ϋf�!�/� Ks��yA��W�/.���@�-X㙄�t����H]�~%��6L�s{<�ǆ]Y��ˢ4�U���묞W3Y�0Ԝ3'R��(�o�t��ڰ�q~��o]ir'g�,���{��8d�M�
V�u��,�
j�z��t�}69�Dv{�d�8#��I.iYU�)�Y��,p�ŧY��m��I�&L&h��B�m��å��T��_�g���`L��kvԠ�tfa��P��&�ӣ��9z��uё��;�?%�o!��9=����IX����}[���++^��
�iZ|�O�QQ���U�����i�k��ʑ�M��� J@^��*�n��
�$¦��͈��c@,ptu|�(��juS)�5�UT�5t��P��_uU#w���²���LG�R����(;�f`;��&��l�����iB`�l�P���K�ϓ�{iN�u��S�ɀ�d_�}��H��=������?����q�R4���l��_�?[l@-��.�����w�N��Yt+��pd�38<��	ko�\֙@�+�>��&�aZ���ܴD����ϚC�b?
.b˶b���ݴ�k1�;�)c 2%�����)RQ�%���oY�W�EG�_�#�4�咬�c������M](U���Xi��E}��1��hdqS����f����k��(��;I�rtM�cԁώ�r�p�֤>?!�$T��9kP�����ފ��jTu��Cig}���M�F�IW�	y�.��j�����-�T�_g�_
���9b��	�j�˅�Nک!��i�-3��Lz�|��H�]��&�\BOZ�8Ў*��FǾ���b:B�e�UAY-��K��jk�k5�7��u9 �#S�1�{g7��	�?�7�-e��ei��ڋ���o!ظ�<���VI�
)2=v�����Y�K`�)��j:(
��m�����Ò?ut�ÌE�x�Cv���$��W��C�s�^O�	�?q��2U���6����{�B��j��O��B�\���l�ܙ�5-��A�䴣�@�R���lz+Kd�A#�S�F~�'�{��3����/ҋN�
�
�״j�ͤ/\#�GwW+���.���ہ����5m��eS�"�f�7���PJ�6~@gi�(�K�H��o�����߭���l86"�-�����xn𘵣9"\�7�P4�:<12��*�(��^SׯF�f���J"�6��-������_�������%��#9|�/��bs/H!%$��)y��IE^=�>�g��C'>�o���s����o5w� �Wga�a�[�j6�:�Ж�9u%'f�D��T�V��*�ʧׄ�b��v};%mp���;���J�Q�w
�����ř7e��9G��Y��	��AIEg����<ݎF<TM�IR�l�uɑ�
���]�c�@r��T��ݜ����Z��O�ZK��&�3��>ܯmJ�j׾�(��� @q�J�5����?�G�~*��D���(�4�2Pi_Q����i�2���E���{���.)ѐ2s��*��S���K-���yԴ�ʹ|ƚWt�rDS��h�=��
j@`:W ��g�FD�`X[ɋI��`�#��p�qFp攩�R)�+��L,PIЭ�<*�R(/镬�M)jh�����,/�tw�F��ue*�����gօ��5}��z`Bܹf�u��S���
����f��I�U�힉��ssSN����/�1hC=(T��+�Y�jyR$���3b��IA��8:����]H���ެu���~2�v��;�����Í��߶k��h�Ŵ*d�{��n��tٮȸ�ZOAo	��4�e���$ґ��:�Πr�{K.��!�ST���� e�5�܅܌��c�:W���	��d#!<�	=���=	vj���|ӁT�i�F��r�]��&�&���O�baJ�..���z�A�;�깵QA��匲�c
���X����ǟ8PT���BU�(NC1Ն�*E�Sp	���v_v��iI�����A(���.-�����ɂ��j�|RR1�]��F��"��ɓ�3H<�7�VKɊ��Y��� um?�����s��h˘�~�t��~v��F�/؀U �ͨg,a?�<+R�c!�\4�J��fz�pN�8u�֡�
�	u0�.�W�Ʈ1t��`�xx�$�7�q�hc$�b�<�%:�K�־�߇󿀷�'�	�u�(�:(���ia���g���c�$`�W�8p�HXE#nB/��R�3�k?�u�m��߸�����-�Z�����G/篫	O1�o[���r9=�N
W��P���cdW%=����E���56�b��`;\3�s�l����5����֌��Ć�Ͼﰌ�.�&5��T�i�Y�n�A�1%�^�^��-�`�-���}-�B��ao���Z4p��:
��'2�|�Son����h����H�ˀrr��)�B�i��r�]&V��R�Ch7�������˲� ��x��lt�Ж�S��ze�E#�3��l�� 3�G��vfQ��PZ�gзC�2 ݑ����.�HM�+��5|D�4M0�*�d�`�B;�RC��A���1��!؁f����vM>)�d����\P)�h6�9��P��2̻��m����h�2j`z	�+�"{n���M�+�3Q��W�]y�R����/ u��2KN�9XLC�*��/��s-d�Ё�?�9���|�1��_te�T;�8Q:�j+���Qu��Ё�d|c�Sj�	]H@킓��b	5m��T�+R#L�����]��7;�<f�f��F#4�$�]��k� �"״cd�(�b�8�8��#Ϳp ҽQX�O"N\�2XH��$*P��EP�c���:]���/T��	�#�q$ HgnDE/6F��jH��{�;�8�.��t��M�^�"���}��e)���/�3Z�7��46�`�����oaIÞ�6��f������5�nwel��ӗn�@�̴) �g2%}S�̬8�����U�j��Uh��lmh�Đ�.�
>=�F�1��9]\���עzB���A�}��I}H��i�ҧy5P�ѵ�+9&1l�.Q�.�|
�S�>=��S�zv�$����/Z�zT,D�� (V�*�ֻ h�M�����l;&�t��J 7��]�'l�H�m,V���M����3,��7�/�Q;�G���F�п�t����W!}�q|�tRt�x���
U��dz�`xP~�;�΂M��n�5��-�'P�]S�bR񟔜�d�|��������
��1��ֶ]��͍�F�4f���C�	Jb�a�E����Q�W�na�~���~�C҂�O�')N��'O|��:Cy=�LY�-F�+�'W�߷8ދ�7�Hn��)��&!�m6g~� vÔ�`aN��뱞	�C��J�����ӵ�{"Y��V�Y�����/�B�/����� �,�G���U�z�Ŧ�dod���V�GutH�⿦!X��M:P��Hk�b��Y����hkﺒ��[��z]�棬p{F��C!��t�q6}Y�VQ:�e\�Z0�TֶRu�C7�1,�b������p�:͡�5��Hɳ�\.
A��s<�u�ڨ ����]ûx����K�"�e*ů53k���c��Hį���L�\�j�w���N<
�����3=��Lusر��2<!��s��rϥ�*�gۨ����lRѱ��1���0�	eQ��/v��%�\'���-�%�w`�����WT�(r��(��B\�~��s�R0t��M���7
��&�w�_G��/u4�u^��t	�����hM��S��i���^}Ξ��S�7`���n��w�!/4S�ܥ>��������0W`� ��w.8���e����}�x%�y��
,�s_�����w�Pz>>����Ot)ìTמy��>6���OS���rR	���P@����ߠ�1(I�/��{3�����;E�f�OH-𧤚��P�������,�ʚ~�m|��)oH�\�QcWO|�ز>��/�2H�����O��Sg�럦��1�	m��m�m<H}��N0B�����^���2�ц��� ЌNu�Ra�[Xk�e s{�x��8&�U�%c��X�Kt�r�������F;kCN1����w����Aj�ɷ�f!LER(�C�P��)!�������_ f�k�����i��+]n��¡Wq.���+n��j�/k��a
�Ew�,���8�� �k[�کӲ,���e�=8� ��CL�4۳v��W�Y�b�b���u��I��$�hw�����_���x�е� �[����#��S�����
��?���\��0��q�*�Aa�>L5F&�Υ|�Ͻ�r��Yw�&% ��@I��
�R���|e��&��mf���*�h�R�!|1*����5S�2�y���np��J1���M�(���!��� (�ߧ1�0���7��X�m�r�"%9"A]P~W�ʧ���5X��ƭ���x$́��T`�Z6�d%������� ���x�D�`��`�iW�a�\MmwU� G\zk�Au��F���o�� $�;��{� '��.E�C�7_ynω����׃mi>\FU�cj��S�o[���:P��5���b�u���;�M�ͪ奒dp��m�̓��[>A2l�I���G���ˎ�ช�v���A�P2��D��a�u]�?���r�!�6���f��ɉ��Y߭��%A/u#�G�wɎ����N���G��ܻ{n- (낎�/�X<R<	�"���8(/�?>C�J��*�99l�E������}�E�2�v�Iy4�2��j�rX�Q0���9��|ə�s5�6j;���T�=�:,�G�\*�f���C+N�!O5Or�<Q�J�8*P�k�l�ʦ>�5�=��O��FU�i]���i#�B�ȣ40P���6�س�Y1���dO�O�4h�B�'TsT�)��B0��d��p�
��f�*|�I S�w��u6��^��࿥i����`�@� �X�N�).�X�'*7�#p������ �����e����1�������J��
B���
g{���">�5������1��Zk��ͦ�	��$T=>������㱴s)�~�R\�����[y�P����T���54��(�б���L����׷���jؿOP��L���Գ����U���!��]bxnP�7��,�Lԇ(�Ta��u:��\C?����b�?�i��q�l��_��s��7�b� ��I�~@��0���(9���$�����PV��Q�]F,ޛđx��H�bB�9-��7�xꄛo��<��\N5e����B��yx)�R����#'6n(U��Tbɋ~����H����P�����F�8	��ւZ�e*dywũύ�mq!@��p���sB�pj8*�����'"�Ά��NV��z_�G�ya�qD��9�<l@�$�  ��v���
���
�	��~I��Z�S��S�5�ٳ��Pd�5P�ow��~`�g*e��y�3e n��e�Z�F�5<�M��:Ns��k9�[�v�i�/p���D��_��4_	{��zE���B�<�,���X�;9D���L�l�'����DD�f��/.��8Y��rڽA���cr`�0�{:5�4ˣ~��� F�Nk�\��tt�ah���Ֆ�`F�6A]�xgB�C]�S`c��H�������$��ۂ����5�`��?�kMޛ9Jg|2���J�c~ð���]��Ԕ��2A��w�~_���Y���1;����-�e� "\n�%�c��10t:��Aw��&�o-���j�KLUl xʀ�����,������@���S��Ϫ����n�Ԥ%ԑQ���M&'a��f��:����������b�|����A��Z�JW_z%j���) �p�>M���c��ທ�6�[��f�7T��n��fH�h�O8f��=���P֠$T���$H�SyZ���&���ݦՃ�뗚O͟\ԋ�з�?C�[�[�BO
^���I��^?3@s�qo��]ʘ��JsY��O�;5��/$s��v����W!�U�sRv-�=�P��0��ca�B�^���Y01�8t���b%��󴷸r�w�Չ����_ �g�J�Ծl����~�ڤ�՛�k������[��>�K7��7�/�x�ݓ���z;��ΧO=瞯V"Z�Qz�6}���*�'Ľ6f?��G �x�W����Ii,\N#m�����g׽��1�\��@z��>q���Q:��� 鷶�������![P�d,ҕ�t��@o���d0�k-������M������FB���[�ʾ��Ћ� ���Ơ�=ۙq3���p�V���1���[��f��}y�e*��T��"�p���vK[i��D�M��5��]��׷W�R?�m��w��6��������.������ݒ̤٦�	ܮ�h���C��n#B���� ��C�UUx��k��M�i"lӵE�rP@`4�6VL�!����-~F�,�������;��&��:zS���<�|�t�ɯ1э��8���r�ԫLCԕ�+���?o$2 L�If8MpB�����mV�{0��[Nہ�|{���xh;�,?�qaK��rJ�x��.����@b���Z?܀%��0���=�h#��T�_��i ��}�
��f�&�R��T�VBV�8Vi���E��[ZV��KJ�wEpKAQ���G1����k���QU l�Sҭ��*�Q�>:�3����;{�\�]�i�v�	���4���u ��T��L���>!��E��x	���%���3_�.�L���^�|���O���S����%��?{S6n^����@gw;֝1�R�]͐M:
O4ܤ����ˈ��#s��D���?��v�m�i_�OS�_]h]��i�y�1��M���,S8"�^�r����M9V���gn��1W"n�rH�뉦���U�R������2�B�2���fX\�N��T�@6��v�2E����#�I��]PGB��_g�P�I$&;^�|.<��M�^�e�E�*ޗl@hތݭ�%Q�Cg�	�=M��$ǈ�ڨ{�D�Gj۴�H����")>��kD�k}�[}�3�,?[h?|n������;����]-
� �� O�c���?^� �������M �aO|@nazM��f~knMN��8��ذ�:.����<]�A�a���ˀI��C�s���`DJ����,����	���N��c�c�u�%��oD�B���d���q�!ky($#�f�5�J���*�{���U.�:���(��+, L�6�J�;�yPn����v��栳�I���n�$5+~�D�674-�?�~�*I��u��|,����}��.~�JL��y�ޠ"f�&��#�D�����L}; ���<˿E�c��W��J�4�d@5��Z�����>��X��/ٹ��b��C�#B�s��1u�)�
�d�t��Ê|���ȹ��e�f��٧ƠE��
8�RT�hf�� ��䵰�$�����sk��6�bsD��~8�����~�X���{��s:8]9j�C"F������؞g��b2U{��'N�oޝx�D���`�}s�	�;�ƎA�PD:�4��v!^�\�	;�_�W߰��h�m�T�T~��1�^L��+w���}|�\���!�(�m9ҭ:Va��Sd��,		XC���J՘���>{!;LA�t4P�d�u9� ^>ī`���~eƖ78)�,o��E[Ia�`3�諊H�v���:��@�r�Xbm�/�.��?�" 6G�p ��ɴ�}~��×�Je�3,o��c��hdӾ挮����#M��7��&�'��Z��*�����4�{$�B{�F�pW�M�n�����+Q���������Ի�Y�+_}8��I�A���E�>�7a�����vL���cS�f��~�� �]�:!�l��W�;ޅ�����I��� ��<?MGTf"��jd���s�T�(�$O���ǭܨ�)^ ��S^��8�z<��I��Mf�f"I���Ľp{����o�d�f���v��m��`�T��q���c���n$IqU�v�u�p�+���dR[��BS�u>5gҳ��ϰ�韢C��O�j�p�TB�;��>�$F�O�L��X�N��"�`�yi{�k��J��p�v$eOSc_�������補������ht裖��0򽻛�aN�?����v�ض��e�мx%�S�d����8��`����f�-��F�������B!î����pLfo�B�1Ɠ��Ea�m��y+�!���?�v�b�H�8p[4����y=J��
�+�/i���<��	Iqӵ�Q�^ʵ�Ġ\�0��U<����-5�H���Utk���>�z�d[D��kc@�A�>'��+�a=�#�A�4��xg���^�@��Mc�I�]��(T%Z?87������I*ج���Kl�e��q�d�����m��E�L��1�"	����6x���&�5�'�D��!���q:+-�нv��ej����!�3�\fe�_UR��"M�G;������c�������Ai���WӨ�� P��oD��˽r�x��+��)bc9�*&�"
( ��hG��^�sO�'s0��jn�0G�Ib	C?I�ՐV��XP�geR7A�8���*5��\�Y�}h� �~R��z���RH��C뭉�Qc�vT*��&6���7{�?�LQ�L�����?6Qj�gL摤�א�Q��^��[o�(����Z@�Xa~[+�),� ���nh�(E�����kewB/.t#j���N���Z���~�6ź`��y�SR��RCk���No�����!��MF�����|]����c��)�ְ�0Q<��vE(��*'�s,���`��w��� �yLo�q�<�X��;���˪Tk!G"Ә���@�Ֆ�kw���_�>�Ĳ�P�ǧ'$9d[&���h.�v;����*{�N6J�j��/;"�����պ���(���F&Q��~���=x��%�4��p��M�љ�yL��m���w:L��A�D�4^��t�~HR��c��dhۖk����=}2�s���{BD~-+ey�Y����}d�����>8A��j�4?f$kv탙�S���`����̶����v��ؾ�̈;I�p7����0!�Z>�4�����R�� �v4w��F>�����Cy�˩]��E�Zؕ���<��cX:P���2%;w�Q6��&�F�]3��SӱJ�ƀ䈚N��?�(-pB3��h���O��]8��Q�&�QI�.�?`��Q�����x��������%�Z�@�%bϨ��u��L�&�) �O��}iۥm&N�(3��\�yؒjdZ�Ϫ�� ˯������T��kX*�Le9��b��rM�������Qq�;�f��浽^#�nx6����F5H2�|aq��b�6Z���k�<b���PaM�v��~m9�=$m��� �s^�'�!��C�`��!3_]��FP��5M���&�ҝ" �=b?��!�`b�u;�ޱ7�<{�"��%�Z��#��oOu����QmX��V��yƷ�8EQR��:\�T��|��g�H�Ow3Y�����z�����0��TP6�T}�{�љ&���s�_��Uk�9�n�L.4���Ԙ�g�s8y�m�+�*�ax޼5 �[��ZF_��.Z8YJt�&������a��vݡ�vI��ɖ[M?(����LEH�p�څnοFwZ 4\�#v�&��W���xrl�a;�h�U�WAb���H�%(��ĆJIx65c�d�
��_ǹ�*WQ�P����ƛ^�N��U�n�u���1F�I�Bzd�s�b��
�c�乙su���V�͙���b_��`�P����]	=<���Ɍߛ���VUJ-��:Q��k��(�㗰��9��ڕΌ������t�S�0����E��`�9*%�-��3
�f��%r�;�����!N�:�b�4e�r�d�$|�w+E�a�~��]2j�rO(_͛�D!�&���hy��k�?:b��;�"��L�R���#�9��s �;�+C���w���u�v�I)z�-m6	�s'�!��k��;\D�e�i	p�ڟ�
˲����SZ�=L��fo��̶��A�m�D�g)C" gEi)�#�rt��#���]��W@�S�VP�Rue~q�]��i( ����5��ۚ��;w^���}��_��-��Kloy��Y�'���V�5yhO����yX�Xd����!�a0G�w����H%p��a�Eo�;�"�yλ1Z�=���0�j�Ȗ�Y;;�)j�蝣M�=A��\���Y�E�s��żL�������0���dt�4
i�����ؔ@-�ym�FW���G/�9܁��&ڦv��$�-�k�p�I�
if ����ucB�W�U�^�d8��(Eb[�y�^j Gs�f��>��N�8=��0�|�Z�8�H��8��E?Y3�{����[N-ZHΡ/d����0�ث0t�Di���5�}��D1k�?a�7f��A��53�����Wnl~�ʧDl�Y~^8D(���r#����8&���@%�^�Df^�q����a?�k�#C�^\��~WP�i;�Z�+��38 ��Ie&>��9�)�B\d���2ɬؤ��X������3�j9����L^&Wm>vX��~�и�N�y=����BJ�>�_�*�0��P�ߋN�,��i/�\ה^�*Bz�����P7k}�b�Ls3�~�����i�N���pj2-���q�Q'��\�����~���Ȏ!,�sK�OK1��L�{B��`������\L�	NU�:h��A���W���dކ�?h���\i����h=#����]#'VX�j#}��p�a`X5�۵��/N���(餦\�ͳ���C����x����t��$�}��Z�̒#��U�]@,7�gy��@����>�5Zg��(��X���p�1��m:�Z�����A���ǌ�����7�C8*9���o�/cł�o�-�+k���qb��-��|N7��t��l�o�.���(D(0�Ɏc�.�g"�»�3lWgT��};�,�v��(�{�4z�:��0�n:��nUbbނ`��g{ڪ�g��4q��_���G�@'1��Ky�^��O����;9��y���������vuڙEy:ed�P��%��%�;f��S�R̺�G*�_���)gH���N�Ϸ�3M����Ձ��aG�u�p\�i��Q��+I�AT�ZtSk��o�����W��v���� �9��[���d�'"�4���k���������_L���!�qcH�c����ĝ"�{p��	�[�#`3���1�D�!�s�k��Okg<k�!��"�Ɓd���M�|mw�|��_�j�Y�BaBʹհb�ޣ�L͏/�4)-�<2�E隆�,�8������z��i��)�"W�>
E"qݸ�9hz�RS�I&"v��'ջY���93*�l.��ј2y�4�e�mu��'�s<�Cd���*��tD�R����%�i��Z��?��,>EPB�BtO����, 8u���9u7CR�����w2�����a�ޛ�pwJ�,JE���>`������(��w�8���,��Q��?�P��$�au�y�5WTuɝ�t�UZ�T٪��u��(�O�s�ʊ#�����}��e�M��S�-���+�f��������O����i�3���L��?d9����X�/\��C��������eVi�Ƞ@��$G�db�#��KQ>�:��x�y5r���L�X��{Lؼ븈���o��2��ԢO0G��\�T�a	b���ɢ�+G��#UK��	��σ!�����ZZ��]_LrΧ�����J���ڄ�E!G�]���؄GA���)9��!��\���H�>V>N����TN��뢚K#'�Љ,Qs���OF��3��?�+Ss�]b��vPW�A���r��(I�5�{�5�)'C�󆇚S(y���2��;�H.�'�W��l��Yd����a*BzdsU�f���AZQ�J#�lW�K<������0�*���*̆r��iw���k��aW�=��ݢ[(������祿PC�Eeg:Z-�c��--/��{h;�\*���DPs�ؙS����~�M��W��Sk	�4%X��/�ª�d��b���O�z$M Q�j5x��z��_{�q*G��>Eeo�wm����}���F��`D��;Chվ��y�:���cJ�N^L��r��ȯ3�o��^��m�]"����%�$�t/6�ج@N�|��ؘ5�|oRl��_��E(J�k�^�2,���P�1�F�������F=��:�}�� ��3'o��6���E��ʜ��ڏ�jx������G5gG��
v?b��72����`x�����#M�a�T�0���_N@_�q�B�o���s{�>�a}�ω���I/R�n�w�˹���=k�C��%i�9R�uy|�/Dv
V���:nt]{]Gq��v.��Vʗl3^��sSA^]� ��ʠhD>���赇��{l�;r�?28���۰�����ı�LǇ��vs uL,���AL�k-{��Fh�l�����^�#�N����H�a�r�쎿{1��o���x���%�ыl�o>�ϵ���"���FQ���
���d�?Y�f�8E-�Z^u#P�c�������T���cH��X���2m0Į��2����,>j�#�?Z����H��Y�.:�הfH�����T9��oPZ%TjU�V��Z=�ZYL"t�x�3���]w�Mŀ�2����S��AғΛȞ��W���P�;�6�����;��ጏ-�i4��n,;�eƕ��a� ����>=�u��x�D~����E\c:}�����r�Y��(Ύ�P���ȼc-:�[ f�"+�ԵF����d9�&ߑ�p�
��G��]�1����ua���!M��d�d&vU(�fd�![��^��B�k�%Tݱo�gYe�pN3v�{��0�˜�>�E��J�g��(?�_g��O�Gʛ1/�)��s=�~蘏���\��A��ާd�1=<�*CMl���W�~����@R�S�T��B:i#�I����u�c�0��e�e�[!�(�6�k滠��(�&���L���7�h�"C$d��Z�"�Dߧ1o��V���$����nlw�u�m�t*�H,�j�TunB�_�&�E3a����[�A��I��>��P+�v�p�im��gO�G��~���`6�\m1(O�E⒩���稢�r|�:���}{��Rn��@^�Ʉ.�e���M5#����g�����8|Sr� 3?���W�H�-��_��m��ѸQ�kD�L3���S.W���Ȑ����(���P�U���fc�5�yzE�
��儁�5>���r�]	~YA������~��"�f����E�u#��&�V!��i�_xF�d�@�	�/l}dW��U�G�/��2/����]n���6�];6�J����d,ݻI?�;j1��8\��+��b��;����{6%���l�#4V����_A\��W�O�����*)�(���D_�BУ��2@!�`��`���B��L�q�L�&�S��A5P6� ���1���C�%´���ܢ����ǧQz`ʣ�V��zYI�-�:��?x�e�2�C�Ӥ���x��7��c�'�b�(��S���>M��CkG�]-u2I9%<� 澤�U`H��%[�~!	�/��-QGD4�T�O~տj�����1p��3���5K�o�2_��I{4�������9o�-��Wt�yp�3ۀ+���g��a� �4�W*	���xr_��dnBQ�r�	e���jnWq��'��׆�,�v�SjcM��l  m͟�)��Թ��YZ�h�S���r���S�������w(J��gH��|}Fߣ ��%o��ы3�x#ީ�t4���3�Vů��E��{�ˎ����~u����B\�v�s�4����pR�2�KX�U�X���@��v�	#��C���a����]�)W�ە9�<r��`�J�3�&b��x� +�Os�~3�#3S��"|�8OY.��!�
F[j�x��-����Q�T��h�Fk�-��c�>W�m��Q����B](Q�U���Q��p�p���PR����ww*cN�N��������,Y��m	$B%!Ԟ 
�bO9c�t�o���m�.�&2Ծ�;ڇ01]��!O�c;���Ȭ^��w�yAm$1\>���_��ټ��Qk�[fc���'۬يD����:?�m�F�|��zF�sP�0��b������IL�,���ϩB�&8�ٴ�z��w��F�˳�2�F���=���B��'��6������1}5�/��J/&,-pÎy�����y�!]nX8���]#��0�$ů����ҟMڂ��K�M�KVH���؅�ަPF��o	�ٵ���\	3-���'@̓''��r
��oB�ۻ����?�9y��^$��26��g���Ym���E�����јN��k�_!X	sv~�+#uA�H��}�������.�Rh�ܖ�^�Zka��(�&hZ���j�8����OcSWo�ʵ�S��L��'_!�`SppE��$���\���l�"���[�A�����O��(��|c���C��8c+�Gjf�D%�e��n�_�2+�u�R���y�I����˴�������3��c �Uc�ãl��@>\S�襊I3 Δ��kg�٦nN'H�N��[� '���J9�f�U��	k�|�Na�iVQg���<��vF��	�sn�5Vݴ�!�am]}�սb�C�w�)�,�M���
���_�E/6f�T��������h��a֞;S��oya�aOCe"6�T���YkG(
l�瑋bgˈ���F����Ŏ7zˁ��@#^wx���vr��ي(���6By�|� ����Z5>>D(�|7�WPu�; .q®����]��u�b-� ʶ�/���X�v�����a�����e���btB��	�;��Td1 O�rս�3���* ��נ����z��W�>���,�O��BW��0��x�k�����g_������A�c�d����E�����l��cz
��l�)��4\�k@�nl"��^C1�W! q���h ��͙�RL�j����
��!�*�?���ldM<��:�;��c��.�O��e��qK�r�-!��r������ �̌��34K�0l��`a"Bh��X�_ݴ.��Eܖ�����\�����7�P��S��$�,QU�Os�U�\���t ���a���:{��*2�͙�i�^��1`7��2ۥ@���
L��l��XU̴�]D��?cC�d->��F��� �w([��ED�JX�x$�O���N�e-wO�7�YO��?�|������*)M��	�dfA�	�B�e�6f��;e�׾���W�7O��+x(����2�V��*�:�i�Ë�����4BX�Mg�O�ֈ"̅_B�R�� v��!"7�������z{m�r�� �����d<��3��|��B]���9�ax�bV�P�S8ȗ����t�|��f.������ʡ!'|�_��͡W_;9$�E���*E�Z_\Mb��O4o�����!\5 Cr�90%���'�$��AA{�|[�ߘO�]�x0At�r�\�vnr����3�
ƫF*���D�����%�����qp�
�	��$M�;�x������3]�F37%�"h���U+�ՀN�˘���e��
oގ"Z�b�B���GmK�...�p�&����+2��G)`�\�j�f�Z�p��=�E��dX\��W;N���"߅����"	�a�UT=ԥ)y�F�^X��Ȑ��z	�����`P��:���y�����x����n��h�����9�����M��|6I�鍐��;ҷ'tM7ń��������zj�w-��hԐR0���.��L���~����m�k�����@x�.����i�z7L�w�8;���%����[Ev�SϘV
0U�,L�~¨�ɺ�)�BX�K[��zC�4�R���H,��Ϡ �!��˧����jI�̳�(� ��JZH�j���`�U�x�WL�ۧ����4t�N�7���ȕ����=[K<�}��8����5�#�5t��8�0��S(媶Q�O[��$��UE�a�;�	0\yXb��,b� �^��R�K����\��UwY�MGn����B���></L��GY���h{��߷"a��&���u��:�ـ?ǆ�G�'L?�o|Q��Q9�`A���h~�+�%�?\��B�d��[���o>[��h_���-)҇��0 �g���I`=!	S$�n�Ч��ǡs gv�Q�m}��`���b����%�<'��O=cVYjW�}؇k�nƿZk(��/[*ԃ����^�Q���Z�+O�y��v;����l����B?f"�ןwR��E:�L	� `�=������i�!�e	��v��Lp���+��)Ų�:�&���I���0ܢi:�9�/9p��&~���ST`�z�t�[�d;C���-�2���2��cf:ptE�L�V�*�T��G]�'E^:��``c��#@�<�����8\Q��Ί�r!�bf`�9��q��w�K'>�k*
�t���=̯|W�6�35�*O�z�P��"-0�G�2��!<�Q��Dh��PH���6<�إT��SN7�ۃ��zɓq���������^�l�fA~N�>1hp�ru����U�3sx��i�$lV,&�S)����n�Z
�{�=V푛*���[�)xk-�u�U(x�H���G�ô�����#��L�_y���֦ʞS[.��5֋��[�K��S�m˦���Y�:ӱ�q��nسs�5��o��b�r����Y���i���tM��9���q�%&ݻ�dQ-o��5f���Y�[�gg�����v'����"���m����˽!��xDD{�j|Ai�m�7���	0���E�f�{�3c�NrQA�Z���c�VC�p�L�նOC���
i�$��Z��'f=��KwrG>��~��L�os�VV��!�x���ݽ��CC�V=�=���H.�=]d���F=D�L9��˗Ӌ��_���	1ihn_�2�Jtp_�٩�$-�l�s#�o*���TzD��x����]Q�����x�����y��8���l�IhgWMI�9��!���p��[~?��/HYiq��N��U--�zs����F�7n���t�������B�H)�k���7�C���[��J��ެ����_pT�D�p�t;�q��(��/U��#H��\4�6�ſ��r���Z������/4�����C��	`A�"�v,q۩5��
��Ut�F�~@_�3a[dG+�(�Ҧ������ ����-f�z1�!��P���ڹړ��lV ACM5׃.��Y<�7���:Q�YAX��Ξ�R�O��i�ܵ���EN��#�m�{\'ݧ���%y������]�~l2v�y)`z��Q�K�(�҆L#R�%�)P OMX�t�_.��L?0���<+�B*�.����a�3���m�?1wW��L#��E��gU�H�'�:�Z�D������m
�l>f�*���m�(>� �f���Jl��!�(�#��43��LVaK�0Ώ��}3�R�����N�j3[e�����jH�Z��tJm93��,XN 56��t2L���bF�n�V���3@"�K��z�[�R<�^����0~.�SlU�Vϗw�E�@�@Y~Q��� �����fڦjs�c4���C��f�9�?V�}�ܒș�|0��	:�@�O���@$��_��ͪ�-a��[*�~Di,�t�P
j��,�s=��ի���8�׵����I�G�l�/��.��'6��������I"8���ֽ�����-��Q�k�)��R���#��Ue9���}goK�d�2ۺ)��[8X���3�����aXP�u(����,u�l��Dpnk�L&����@*
#CM^���U#�?�E V$'@�;QQ�D�����_
�"M������k�w섖�(����W�E�l3�θU�@L���,��2Diu}F�S�.1��\��x\�����{v/S�m�.��%i��;WIQ�H0���s'��gӓ-f�h���.ᑻ~��J2���`#�[��uXr�:�}D�U��7�-���K(��clo\z�a|�x�^�@�s�gE�>~jf����{ ��c���F%~�i%�-������H�L�����{e��kJhlio�ߟ�AS�-~����!2��o��Ѡ���Y�W�	�B��Ӷ�?{�,�r����}�$�>"Q������`�eo�h�b���w��t�@V�B��t{���&�b�t<Y�N3�^P�m٭�Wq��E��m���eՃ|���|6��ov|Y쐛�v�+'��x�<����B	�Z(��W0�Yv���������'-l�P��x�x2�����~�ʜ���]=�|x�B� �7�>K�y�/�ى6�N��f�u{��-RrZ%T5}�f#a���3�K�:H�Tdl��р�8�
D�J�|�����p#�i�Sj�/-���0u��kRcf�"���J����}
�s�E�-Mfn��k~&���7���}biŅ�O[�V	9fu����"�-Tr���o���Y�?'}_�����~�3�j 􁫴������C^O�H�mc^�{����⁁��T�h���4L�.���* �P"e�8ɵ�a%V�P��`�p�� �f�M��
�h��:�� �9����C$Q%qd�F�O��Yp�ep}�vM���1���bT�o��&�/�����e�K�x��S�$��r���gb����[���
�b�ֿh�T��n6�Ը���S����B9�I���"
A��[y�'ڼ*��(�'(�
;]6���	M	?-�����>G��ت�0Oioէ�X��
 	]Mr��1��ڝJ�b<Z��!b�l:DE�u<��4|dK #�����.K�F�z���Ǜ�ɤ19�?Y����y��niO�7�Z�Dm*D�� �32g�h��5x�� #�WMo����
�hq\��x�U^��z�C�M���gd�ot7�X1���a?)n��-jj�����J��lD�څ�Y�#��U�W�XR�7�DN4m�'G8��,���/}m�0f�#2Cw:I��8�$���|
q�	6i��� ;���}�/�qRɍ������=�d�z�3�5��]�'���R_Դ�+�=g��e�G-K���]�|єm��-Hi����"�$v�uA��K'e��� �EK.is�M"N쑁��<4(�M�+�=hp8<'g�a4�Q+ۙ���R.��jױ�S$�GU�o�'[96�Y}�Qn���\:�)ud-I �6��nc Lqda��n��y	HÊI��h�'��7V?��B7G���ޚ��n ��IctpZ�g���V�e*�5V���-��+��g�� �OHt��Y�zA�rx��Y�_K��.��hb-��_�+�l�╂c����t�Pql2L�e�ߎ�qv�t�=:�����Y�}�n�Q�8M �芽�}L�i)
�C�|"������_x��ٜ�q��]8ju��%V��fW���) �l ���4����^��0T���3�?A֟�G����k�?����&�w�Y�j�����
���nȠG�{|�a0�V�l�c@y<g��̳�%�~�w�;�1e����#S��暳�p&<�\�$>�T[b�9N*�%���z�;�`�T6O p#��%�\�K�L�$�a�6��R̂>���:�N姶��^g�r�c�eZ�A��?���(�?	��[�|)�#������(w=4Ό^C�K��+J�X��B\��������k�2{݁���y���q l��h��@FvU����EԈ]�AT� r�K�1���a!��"��/�~�-mOCY��+F$�O���_a8��Y&�
E��ӗ��A21�*"\s�L�J�St��5���M'(��xY�����g'.U�2{���K��������O�H� ��umz���f��b3�����&s�!vO�\<�S��^�ċ��y��Y�!�%���lc1ev�Z0��[������T�.sTQ�|�*�{�|�h���߀Õ{�?��#r�E�&��C!�\���^%��b����Y�ٿ+�6�0J-Y�RO�%C�Nѯ�F�n��*"�ѣ-N]��g���>��JO�n���̚����0�#��U���Z!���+�c�'��Qf�~����F����>���Tφ�ۅ�]h��A-d�
!�4��sQ+��p�i��2�F|ǭ��+�������G_�0��M��y���Z�v���P�C�Q�w�9���Νɬ�i��/>q!:���"l"	!'��i�@o/�ς��$اVm�%Mޓ��⨼�b���4h�ީ��n��N#R.�P�%;SC˔+�l}%�����:�/-�|�ҽ�(&�C�M�J�8%2�y���5�RF�ڕ�k'��[oO�4l�*�5S���BW�H��.�j:MLQ���� ��)�F�\`�-@���X�0������Lj�5���ӹ�ݨ�
=Z��f��aVV�~)�,>�!����}GE�?z����?���?�+Ҹ�b����v��7y�sdl�������2IJ��x	�m�	���EGC뼰k'3A�b��-3ɺ�?2��^I�/��c��=^�R��nF�X:�ӼT�kP����)��摾�w���e���m�{
�s8�(�|tsZ흞^h�A�Ӯ��[���m����
%�`<������In�RB!�ͭ����p]�g[X����T�M�_�7*��1;)H�R ���yf:7-�S��J�>�@ A��AW�(��٬�_��+���8s��,Qv4���Ҏ.���uX��%s�5������/�r ���<��`a��İ��&x�җ�A l�O�d��9�6�EQy����,^�̃�|�����9&��ށk� Kƽ0ÏQ��X�p�g���%8;{]���qIO*Z?��E��%�ΰ�H���+�����x�#.󡭕9�31�{�\�O@�Z��Y�)s��;��ȳ��)ʾ>�i쁋98_i'U��s��{�gv��I퇀D�Nl���Ҋ�ri�^�TAV�o�C�YV(�б�#���,;s�~^̭�����l �[Yɴܫ�]�2*�;�>���P�wLR�N~���=e%�������k�4NDe�m2�
k�y~�,���dx,`Yy�x&�׫T����$��ᴄ��$�G����|M�w���`(��ͩ��ꤚ��ܳqC)��������ζʵ�3@M�J9kR6B8K��r0���TM���F�-�Xƃ+j���K8m�v1���T����don�E�^�;Xv<�MS<\ƛ�ļƈ@h��Z�l>����~�:Sqi�d|8x����:���wB(�3��=Z����;�Z֫U3�:��}6շ�%�c"ё���`ێ�����G� ��\�i��/.y�=&l"��+ s�_R�H*�hG ��,|O�٘����,����ܳ�I�B
k�ed	�#���nP��M����1�T���.���@
�Q�r� ��<jNZ	���A�քl=`���E۵Zd��u{�dm|���qӯS��Z�y��7�"V�����bRD�+����~e	��*=�L����L�1E��_]�d7��º�%]`��ɖHt�W[�s�P�8t)#N�H8q�$5c���G��|oW��b"*�y�ۑ��/^�����tP�U��r֗�Dl�%"�[*/����M�Q�V�6w��M�SrV���D�+3O��ɞ뎠���#�F9�i�L��5���?��+����A�|��	aSdp��a�P/MJŖP&�n�&� PA=���5�<s�J|��;%\�.�q36jwi
�xЩ����b��΋g�T<Cp���������*�X�Q�,�������6�7�91�$�0��w��7�O���$�r9��>t�O�@��S!���e{\����Z,B�7\-
E�].0OFkbU�E)�����@ٻY377@�a�"ϖ�~=v��O�*�M���O�G��_�h �hP�Iz`�D��]ŝ}�cUj��ۢ���Q��٠f9��21�E4�u���	��Zr}XD�-C`1��^F]�����A�%b��b��W���`�v�V��s�9�n�,���X���ud�|���.����k��|�N��2��Ce|��#��/�<��9x���|�v�?Wp�zٕa^E�!�<����|L���2��t��M%�y-h復L����%��秊_	��Z��g�.x
|��d76�x���c���@o�P&_�Ԗe\�ɬm��4�
�R.�e������zK�N?L�B��J�����~�����?Yy�+��C�eS>�4��]&R=_UX"�Dփ�f�B�:-ʹu���fU�
��_M�c��¨B���_ʨ!x�j�%�ql5�ų8�
�qq�cRt�n#x���Gg�O��'��8��^ [K�{��0��ui)m��Կ�f%�e�ZV���'F�ΧQ���d��ޙ��E3~��0̯��0C���_�[�p�g�򇁎/n
G��AF�L�JY`��0y4��I����e ���Q�r�A�ȑ�,^��G�����!Q��(�w�����,3�G��F'�CT%�ai��#���#�Ǧ䆅!��bB$��NE)ꌿ�:�ZN�e
%�&GB�ff�~�M����1��}����X+�/N�;�����B�t�u�qu��5��)cڪ6�qW[���M�	#�#�)�x&73嚠��#>�a�D&E�]���6�Q�6o�Q�8�6z�37��}�<`���~ �𱗊��5S��d���=IA�A m�}��1���.6�c���ƃ�8Lo���mN���q�gz|U�A�x{.L�T�"�_?��*2�"��=*���i���3 �q��y�<�_dk�������68������g:�������I.�x�1O0u[�
Q�1֖*���
<|�{o�+t�t�qe:E��Q}2͇��b6�*+��,�a�d�4nZ���MC�B����j슪�:Fq������j�,���)<��c��Y~ vG#��I:� ks;��p�[ż�ϳ"��
u����0.<iB��y5�eĆ�P�B�SZ ���O�f���2��x�`��&�+���?�FU^ڃ=�?����X� k��x<0���0YJǞ�����ҘC+Y����e	3��'8㹁���(�M�#��_��`�1X˄]e�S�*u�� �
a"c��*�ڂn�vAk��T��]�)�oϒh�Ru�;��|!���~�������r����� �X��H�{����	�'�_�XB��&�:���\~�O\�QE7?��=�q=�)׶���)�Ad�:�lGs��9Z��i[3Vߐ�?P2��� �7ohv@U���3ַx�p�g�kh�:6�Ɲ�g�0�f�ɦ^Ʒ��8���eאyWr�p�4!hF�§�L��N��	�T���n}�٤;D``��w�!��A��_+:s��i�������#Ԡ?��r?<�м�k+�8__���/^��`�s�p�b�������Q��P�C����Z�+g۽¦��m��n7Ӧ�J:9<{���F3 �r���ǒ��ǁ��������)�`�<3��Qֵ�M�0Y��O��1Emt��c�[ӤP��b݆#*��on{x��	�)z8��f;�kģ0t�3Ü/��o%�auI�m\��:]	��e���4�N�)ΐ��".Kt�>�A�*�� ������↎����D��7��%T�U�X�_��x��	O��e��j`12���OOř�+!�[�"�m(�)�J��7RQ���,�N���������wŴ�����c���e���`	e��#@LʬG�� �����0����L(��ňw��yĚd��C8�M䘘g�|�k~H._��$Kh���:�G<����,�
]�n�tp���&_#���s��v<]z$���2��v��)�Im���41�#����#�5OG?$U?[G�af�齯�A���(�a�\�l� ��};%��i�1�z%��h�r{81��q�æ~�r.jU��kvT4ݘg*�x�G2��\�A��M�	�,��G��)X�^=�#Z���wZ����"%������)�|��L��L)�1+E�;��0M�|A�w�_R$�C�G
q��۽3	���
ɐ�<Y.�~�'��n�q ���Nʶ �b���`>m�@��p+`�N}<���C.�駍���l��D�*B�ȑ�����r���h����/!��Į� ��a���$��.��!Ұ��B�n��S�GԞ�++�Xx�b���z֚X��?���a��%���[�J��A��,S��`g�:KW�s<߉K0�B+O�m�X�:��=j��䝨n��D�l/�Z�u*(���j�����&F`݋�N{d�4!T����@�H����޵~�>Ư�����:�J�
�+�6ſ������������n�\�#E��f�{|62�D���]ѻc5+����i��;�Fyٱ��,b�&8�
"������ĩ����߆�G?�t_"j���F��G��:.��"�-o'@4,��,�ܘQ�A�{"/Xk����-���i��b����I�HR� ĕw��_U�tl.�f[W�l	x bgP�9g��t��[KMI)e�p�3$�����¦ɍz���6�.(+�UD|O)�N���ҩ����^>|9�:
3K)ɴT���Ki6� ���G��BF�c${E��:HR��^�VEV��S�rڲ^�,�
1�*�&B�٘YJ��s/���y���(s�ebn�� ����P r��4�����w��� �.�?�.	݃�).
�哎�5M�~��:�b69һX���=�\�J��2#�)Qw�>_ �� ���W�z����TI���VlT�t�:X�j�9�Y3]��濨0�z?ۄ�\�u�+�'ol}���$���cEF�K��C{)���!kQ�;�2��+v=$���&�ka�d�����t�B��m?��IG��6�b
�MoJw9���pAk�-๶ޥp���ѝ��Cz�8��Beɇ�H�r�V�^��W� .�cc0�HQX��4ӳ;��(�7� ����E*4�^k3+>C�xj��C<���5�z�0�\��]B[�'����~�nEl9�z�^2�:��ŗFU�S�c�&p�o�w�ː�ׇ��H����g�A؊�;��Ѡ$�%��)�M�	��"�'��j PmoW�ls���%]i��7VWP~�z���|�DȻ�����&7��m�u�X�??,�5}�2�������:%8������������%����S�af�$?��)ؚ.m<n�
g��e/ɽT�=�v�z�?.���n�mB���Q��s#{|&B�bT b��4��=a��,�Τ���������sa;��w�j�O���(И�B}}0J�L�����
9�{!5i���k������e[F5ٯ[�7z�&�z��$%�!AQ|I�8J�"��)�-��j���GY<<���1h��=��Cl�h�A�RK)���2}�`x;,�	�uf�<�{�}�~X�,u�7�{��@��.N��x�705�����)W�)y�Iӻ��b �����:H</��H���j��hc�
/z ���rKQDE�PYZv��~����q&{��^��O�#�h�%�2'�W_oI�l�Qeq�+*�2�"�=���c�©{���ʮ/�4*��`��Ob}.� 0�t���ٽ�lX��[�c���W8�W+W��UЃkL�����ٙ�~�Ȑ������I�5� ��id���д�Vw0��;F��S}J����W�@��J[J�m�����O9��6� �]��&���ɱ��Z9,t�K8��,�i�1�$���U���՝��y�o���Fݧep��vWt��x�+K?��XSd0�X�u���[)��i���C�\�DXӍ�pF* �!G�7u��~�"5���@d�_=)�I��k��-W���/�F�K���g�ڱ�S6gQ�%�vӍ@��E�W�s��3J��<T� G��Ԁ���5��ۂw"g��p�gx���t)lS�����kM7��-�.8����H����qhx���|��&��	6&8*�s�#��Յ:������@�M�|((�b�lE�eəv��`_0{���+��,���O��p]�8I� ���
��*�ʋ�ub�(���֕	l�C)�]�ge�GEj�B_�h-���ɡW�W-��? R�����s�S0�����p�Kb��w����T�8�T�����G���,����4D��&h"�s��a��_�I����F�ڟ37�B��S^�ζ��� �?2ե�h�vrBm���.�6��-:���(�����ܖ'�J��8U��_��o�����M�j������Q�CKSS�y#[*�͂��k��Is��O��d�c�c-t?�ҙ>R
���5YC�C�a��v`�T����S��DA��b��ž�&B��!���ю��wjL����,�=�5�tKlK<|�[*e&$/�KaT����k`dz ϛ�䥠Q|ۤ�|����M��?�n}��������y��Lyݣܼ����U.n0�����۷ՓO��O'������3gԉ�r�H �2;�h3�F	�Z(X�|���cR(i}�һ�L{��-W��Ū�V�ц��h=�+"E %�Q��l�fFw΃���xª���ׄ�nJ�F�]���<�R��������ʓy�e9Y~{/�
_�)��T[�i��pA�<� c	<��=hVQ�Dr�~�����Cp#y?S&��՝�a�uM9w0l���v�:��:e.��j�h`��t�3	o<0%^<(m�3N�����0Ԟ�"m�Ԧ�[���KfنBi�A�W�8A)�D�C�V*�ZM�{kf�!c\!P\�"�ɻ6Ժ$Q
�$��2�8��{p;�W*���D�>־���D�ʩ4�QG��rW��YIRto�L��Y 0g�h�N�u��� 8;��7�@��g�1j�>�]����;S,���g�Z�v�����%��ָ~��0.������LQ)�|^�m�)��Ρ��6��.6fxr���9��'��QA&�ڮFe�]�!�lʠ�n�@TK&�o�P$�A�c��c�
�' ��˺�ϧ��?�n�~.�1��TE&�af]�pk(d�'Xf(jT׹��>���\���*����|�� ����K��w���#k��Zl^�j|��}.�51�y��i9�I�����M�о��Q��y�@�"�\��8+b��7��LU�>��r��y��3�1CW�o͠�U��/�(��2r��G�[j��S���Z���WOE�\�w&E?ֻRm1?��8���k$Lf���Z-����Op1�9�(�r��C�2�b�Y����QW�/V����8�� U0� ]'@`�`Y�⵬��+�-�O��>��7*�Ѧ�عE��S��� �ik/��lN�8�I�aօ �?	�|����0�'����5�?%��Z}��t-E"�^A��xw��;D vX��:�d���QR��H�y�[b�� %\��#ճ��S�鄊�_��5��ϧ]��P�X�
|n�aW�q�e3����r�,Q6�	�o�����i�it���F�5���[Zy��^��d�3��a�7n����Ywg�`o�c��g0YkG����۽vʣCsv��O�q���v��R8FQ���U�m41ް x��T74�����0VϪ6yO��Y���6e�ʉ�
�w� O3+@88�7��m> ɵ!c�'���(�u\%�9�����k�����t��}
?�C�P)���N�e��	e��BD�#��<��;�l�/i�ܕ05ح9Ql���Þ?,�v'�|���@�����Pq�Yb&k8�С���Y���e�2�-���hh~��g��8Sq�U�OC�Q$�8�=Q��y��Wգ&���&Y�!�y�-	c^��K�gR��hH���V,ӝs��V@�^7��Bt���n��Awߦu�Ug�u����ŕK�&(as�����>�D�A~��&?=)��͕j#�4��Z��5�M��+vvG]���* _��ׄ~p!�|�EIB֭�6�ԫ��H�G8s��q'@�3*eD��@j�^��_z��d|ӈ`�\���7a�|I�Ų���0H|?y��.��I��(ؐ��I/�0v`�������"tPߏ�4�HޠL��� (Ư��s����ȼ��:�&L�wf��fp�P��	��Ć>�z�X�cx����f|2gf�q �L�F��|`	;��Z� �H&W-q�J�s.�ݡ�6`�<�Mv�ˎ����K�F���U��
���~�[7q�a>A�	��l*_��":�?aٙrc%���>�a���8�����B�|c.�~�q�ח����&�����e�3S��ջx7�f�l�弹����@�|��_
���E.���:)۟dp�� @eK�������VMY�xk:�<�����<�-�}�
��;��VF�j�rdj�Y��/�wj�j+i��86��_{� /F�Eu��/��ѩ<�KEu��w�$5��DO�������NH��P�a�=d��{Z
�? ��E��Eͫ6N5�yW����|��1��y�:��9��_�Ō�ߔ�%�/���`NX`�ܦCP	i����6�A��<a�JΕVy�[,����cSlӚ�t-Uf�Op��O^_@�и1z�VR]w��w_	n�MX���^K�@�=i��S	�|�_?��a�"�
7v�0�R��s�;�ޔ�����VɆ"ú�_�VM�ں����$��!� ���R��L͕ 8�ۮ�ހ�����%�$^�̦�����`&�L�Fן|{Y�N�<qFr��5����|��?�b�G��=�ml�Y�~߾wC���\��@�9M�3p���!��A�]=��N	\8�7�ǇI�B���AU]�w�^ ��gO�][��AY	�$dG�j�~��0$����1)�b��w�:8�Mc-IrZ������s"j[ѳ��[��;�']��M�:�DW�w��L�59�4��o��8�(<��� �S�vw��6�30�<zo�����UTa�!��O��>��K�����J�-�'P��Z�d�^N_�;2V�t��T����{W��w���{ T�����6��A:朗?Ş�����-#x�GM���!���|�!��;r:R6�p�:ʟ
��;��k�t���P�(wv��NB�l=��hgޖ��%_F`��Qr��6#��~�N�e��H��OC:}Sc&�C)!_�Ip���f��?�r���TqfdB��0>Rd�P{F����r�k�>7��6��s��{��e���$�bxΗ��@e�E�y2_��@Q]X�� W���ǈ��W�Q
��a���Z�|H���;��(Ѯ�&A3�D)�*L�<��+�7H�u=y��H��a�Z}ic+L�A��+'�cf;p,�a�{�(�x�h��g�C��i���}2�oO��X!��\{�P�kK�G�T8�֩��j#(�7̞ @�c�&V��6���y#���n���&Ь��ǡ��(�]b�`����c��GGn<Ƒ�˿�K������~�RBE8d�����7	�͜dێ�o������f�n�\����a�	bVx_�W~�Js�la�ٜj��&�`�*�+"��� ��Q��/-9@��-���<ٯ�
�I�!��@��V1#$-/�UID��<�8��l0�@�*=)�K u���%^�d�e��������0s/��]f������.�K�DW��٬�Sj��_+��ܵ{U�����Ɍ0l2'�r�Vf:m pȰ�&�V����{��`KW<)9�_�d_/�!�Q��ĕ���<��q���ƈ����	:����PN��m�N�s/��"q(443A,�fe�q�mYN��t�7p����y-&��+����.��P3�����JnG3�q��5��\�	�7[�f����М��N��R����9H�#ڣ>��	�9`C�R����Y�Z����#�:�����i,kinnW��B�V��0�r�9�3�,xÌ+�P�)8��G:�d�����d��%j�k�z]����	+�I�����~wvx���:�K�>����(�c��8���Li6�QyG�;���.��]6,�ko:���E���VC�N��4��wq�����JN�-�4;�Ax��E����u��8(L��԰�c��ݽ�˓�+�ƌO�-9��t�����͵�@�����
Z�Q,��O*�p��i�����\G�tm�(�|���PF�V����n���qq���v�D!�cqK��d�/�\�Xru��@-T���hi�+��(�c���p�`�;���=��%��ؾ�5d`��m� �ސL@.��P����7\Ǵ��ڏ�,����pJ���v�B�'b��X����oA�	ˬ�u��� �W�Q�yU5�~v�<R��g�������_��b��V����va��H�D{�kK-@q�	�\$$�˗x;uILy:W�%����3)�gN�`S��qI9w����@�d쿊C��g���\�����b���A��#�8�U#�c�FM�v���金���q�,���`���$��X$9M7�����Ǆ�jA�s��B4D��#OP�����Կ�)�)�3e[���*bh�!0�'%*Lb�1�*�MV��&ٛ<سũW�˵��e9L{��W���(]f��l��`�BsK�������rS�R#�AG�a�>9��R������ ����|L>V�fJ���u�:���.�fȥ�/5��;�3�\c�&�H�$�i*tO\S�V�,��Βu'��C�WIZ��Bu���鋪�p��'�Е¦iifgd�y-�$_�y���*=��K[m�\�c�������J�rڨ��:�Jl:{�Eۥ�Kb]�"���ĤN�K~��m���^��d��Ee���o2.'N�fhͤ�WSd�<��hzj�´���3�X&Փd|~W%�5y�z9�`s9qv�mdr�N��r_������Z���������;C�?GMk��/Y����{���izm�.eV�M�In�4Ұk��Z;�<�����gGBO�!���٫/_���;�v<��G��^P,v�o�mqRU�js�8�F~k��w��5Ҵ�_�"��G3�A -,0�����j@�96�UQ�EI�(�}���t��/�ƈ�9�Fx�X�E'�N� ��P�Ϫ��(�6���K�A2��%H`c���4��"[V�M�ʷ�K�+~fr��y��q@�TC&����nzՙ�d�6��fY�R��wͱ7d:oC���ixtܳ%a��l�Qz^U�\��w��,�[�pk.f�3�@sZ�A�_P��}��R���T�Q"�2Z�Ȩ��FG&�����B)v��!��0��%/����~g{�����"��Wmn�IF��GU�z=l�U
G@���(�&\0��:� 2s��[�{�\]\���O �v�ݶ��"�))�Wv�*�ؗ)������[g��],-�xt9J��:�a7{́=GWT}�ȓ���/DpH�����7L�8����H`'�?c��xS���dLS���«N�OT���"č��!��8����K�!�<�U2��Y"<3�
�m������qMR����ާF�� p�()LP����m9��̱�N���L'�0/�FLw�op(l��ʔ��X�_�"+1?i���Wxh^�[�sN�s��nE�p��s�|�W���`1t�F#N���;F�f�_�1��&�Rk�`�̩ ��������\�������e��"���㍱���s���%�e��}���@3��E?��)�վm��&��q�z��H��![����$xe�#�#���tS˭P!����`T�Yl�~�XЌ��ŧ���Y����/~�����T�tag�j�"����TW �Bx�ӌ�"�C}u��}��<v!�������3�e_XZ��}��G���o �m���%���&,O;�c��x�+7R_md\ry+��0�ڦRЩ�c/<�cAO�0>Cv������/}נHq��GS+I��N�����%+��g�j#����J����ΐ>!3��l,p�������w̡`�
�؂���V��S�	��GN�W����[z�#���J�eL X*P�MXl�	�'@���ᇓDeH�F ��nB�d��>MJ	d�c�+�-]�S����o��3J����W2����Φ�a�yt�p��LМ�9��Qq����C������O>��פu'i��jNa�"�I�Y��4�%�|n{�rz��K9ڹ%�ƃ�n"\�y/�"<0�8i�`�KU�S0Az��e�� v�H*��6����7�e|�w �ϛ(H�0J�O�H� �A��ၰ�r}�<m��0On��~����FB�h1���**���r�lAI���^�p�$���	��SӚH�����CP����_��j8#�\R"k����y����<���iuu�w�
��u�X��ɧF��8pWgH�1n�C���SW���
ұ�TI>i'�'1�
JU΂@G$�YK����Q�.Ѓ����>#�F���Up���p�";�����;��6vM��s�5�X�e!b��,�e%�;Ej]%�d`�plF�l��Nm�Z���	�/y�*IF�/%g̬�7���%�a����J��r���m�Z ���G`Dy-�S��}♵��}]v߄ӝx�ş��j��������ٲ�Qlc��dn��`���u\P�axV- �~����Mx� .H��D��٫L\
�r�\�õ�8���.^���y0��z\A��-��/㦵	�H����X�7��[ȗ�bmL�ٕ��r*
V#/�t�k���6$¾��֒� �:+��w��&��иΆxpT(���m	�ܬSo��d&h��9�$ ze2�,����	#�f@�R�"B�J-�Xc�BS���$��!�3$*�3٢N����@����}�[�~�^��
�rB�9�l��rAf�T��S��
��]�Mݼ�2���<�^ϓ�" c�_&[M�H���~��MS/˱�q/�<�9w�E��c�Z'ї�ч�����K<�W �u�����Hj�"&Q,�!Vp�f�S⹥��ͯ4���
���m�������m%^k�{ai��0�������1�y���kr�97��?��фgr�b�;��}����?9�j�������_�G����(�b5qO�?�k+&y�b[7j��?^�%��Gw�(��%8���	���-���{#j�-�?}l2�����/L~7�}_�Y��WceO��^�����v�U.��bB�(�-0s��^!��Ƃf��v��b���ٖ@JrP���x_hj�*�:k㈎�#
e+k7Pꪴ�a�rtz��f����P�Un�3D���h�k�tT�Z�|z�&�(�+.�?FkSbq�i��.�vw#��f����ݚ��g	q⸫��H�˄z�	>R��s.�c��RϢ�l^��Ȥ�̸9,c����	>}�E3-��ivH2�n�V �����!'6��&)�9{��C:�G�\Ct!j#$N=�,��ߕ}��ܳd,�� W����Lҩ����������¥�@ѳp�1���.�a',R-�~0���ۮ
�V�Ԣ�fM碜�s|���r��O�����։^%����bCQ�@4��(�T�<E�v�ҷi$ܺ���)dł�#���_�6��]����ER�>��Ww�g\�g޷�P5L$�k~:%N.vU^t���c�
>�GV�_���Á]�ė,���[PQ aE	)9�������=y.�<���)z6�OP��&��������@.;�-�^I_ڄr����0-��̃½JS6�]��B���� �rv���Ln�bU��!ծp�`����r9[IH�[�_�|�y6%��V������S�2:3�/�^�IE�;0��|��,���q�8�{�'�lzN�B�:�D#sǏ��U�b�P������c\��bR��*�9�~_��T3���ؚ�q���`ՉK��>��-��^�T��e9���Q>Eλ���Z��nF��ߎ�ҫ�aJ;�65����FK=���#m��Qr����s5�'�2���\�v��d��Lj� T��jA5̱48�a*��ړV�yP�%�c���g)���\4=x(�M;���B`�>v�X[�� �.G�@m�
��р�:jJ�ܫ�I�:ںm� `H�W��w���c�G���RSs٨m�@{R�@�����X�&?�ြ��IG6r�^C�c��A���(v��d���
���=���&��lwL^ĴV�;*�q}Y6M��#nK�<*��
;~�>�+��4qw�+RH�m��P�f�D��٦�?J�X8K�tzU�2��&a��CzH)�=�m	�#qM�<�0w���Eox2�'P=�N��